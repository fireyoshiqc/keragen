use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;

library ieee_proposed;
use ieee_proposed.fixed_pkg.all;

library work;
use work.util.all;

entity system is
port(
    clk : in std_logic;
    rst : in std_logic;
    start : in std_logic;
    out_a : out std_logic_vector(119 downto 0)
);
end system;

architecture system of system is

component conv_layer_mc is
generic(
    stride : integer;
    filter_size : integer;
    filter_nb : integer;
    input_size : integer;
    channels : integer;
    dsp_alloc : integer;
    weight_file : string;
    bias_file : string;
    input_int_part : integer;
    input_frac_part : integer;
    weight_int_part : integer;
    weight_frac_part : integer;
    bias_int_part : integer;
    bias_frac_part : integer;
    out_int_part : integer;
    out_frac_part : integer
);
port(
    clk : in std_logic;
    ready : out std_logic;
    done : out std_logic;
    start : in std_logic;
    ack : in std_logic;
    load_done : out std_logic;
    din : in std_logic_vector;
    dout : out std_logic_vector;
    addr : out std_logic_vector;
    out_addr : out std_logic_vector;
    row : out std_logic_vector;
    wren : out std_logic_vector
);
end component;

component bram_pad_interlayer is
generic(
    init_file : string;
    channels : integer;
    channel_width : integer;
    zero_padding : integer;
    layer_size : integer
);
port(
    clk : in std_logic;
    ready : in std_logic;
    done : in std_logic;
    start : out std_logic;
    din : in std_logic_vector;
    dout : out std_logic_vector;
    wr_addr : in std_logic_vector;
    rd_addr : in std_logic_vector;
    row : in std_logic_vector;
    wren : in std_logic_vector
);
end component;

component maxpool_layer_mc is
generic(
    pool_size : integer;
    stride : integer;
    input_size : integer;
    channels : integer
);
port(
    clk : in std_logic;
    ready : out std_logic;
    done : out std_logic;
    start : in std_logic;
    ack : in std_logic;
    load_done : out std_logic;
    din : in std_logic_vector;
    dout : out std_logic_vector;
    addr : out std_logic_vector;
    out_addr : out std_logic_vector;
    row : out std_logic_vector;
    wren : out std_logic_vector
);
end component;

component fc_layer is
generic(
    input_width : integer;
    output_width : integer;
    simd_width : integer;
    input_spec : fixed_spec;
    weight_spec : fixed_spec;
    op_arg_spec : fixed_spec;
    output_spec : fixed_spec;
    n_weights : integer;
    pick_from_ram : boolean;
    weights_filename : string;
    weight_values : reals
);
port(
    clk : in std_logic;
    rst : in std_logic;
    ready : out std_logic;
    done : out std_logic;
    start : in std_logic;
    ack : in std_logic;
    in_a : in std_logic_vector;
    out_a : out std_logic_vector;
    out_offset : out unsigned;
    simd_offset : out std_logic_vector;
    op_argument : out sfixed;
    op_result : in sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;

component conv_to_fc_interlayer is
generic(
    channels : integer;
    channel_width : integer;
    layer_size : integer;
    fc_simd : integer
);
port(
    clk : in std_logic;
    ready : in std_logic;
    done : in std_logic;
    start : out std_logic;
    ack : out std_logic;
    din : in std_logic_vector;
    dout : out std_logic_vector;
    wr_addr : in std_logic_vector;
    rd_addr : in std_logic_vector;
    wren_in : in std_logic_vector
);
end component;

component bias_op is
generic(
    input_spec : fixed_spec;
    bias_spec : fixed_spec;
    biases : reals
);
port(
    input : in sfixed;
    offset : in unsigned;
    output : out sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;

component relu_op is
generic(
    spec : fixed_spec
);
port(
    input : in sfixed;
    output : out sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;

component fc_to_fc_interlayer is
generic(
    width : integer;
    word_size : integer
);
port(
    clk : in std_logic;
    rst : in std_logic;
    ready : in std_logic;
    done : in std_logic;
    start : out std_logic;
    ack : out std_logic;
    previous_a : in std_logic_vector;
    next_a : out std_logic_vector
);
end component;

component sigmoid_op is
generic(
    input_spec : fixed_spec;
    output_spec : fixed_spec;
    step_precision : integer;
    bit_precision : integer
);
port(
    clk : in std_logic;
    input : in sfixed;
    output : out sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;



signal ready_s1 : std_logic;
signal done_s2 : std_logic;
signal start_s3 : std_logic;
signal ack_s4 : std_logic;
signal load_done_s5 : std_logic;
signal din_s6 : std_logic_vector(8 downto 0);
signal dout_s7 : std_logic_vector(79 downto 0);
signal addr_s8 : std_logic_vector(9 downto 0);
signal out_addr_s9 : std_logic_vector(9 downto 0);
signal row_s10 : std_logic_vector(4 downto 0);
signal wren_s11 : std_logic_vector(9 downto 0);


signal ready_s98 : std_logic;
signal done_s99 : std_logic;
signal start_s100 : std_logic;
signal din_s101 : std_logic_vector(8 downto 0);
signal dout_s102 : std_logic_vector(8 downto 0);
signal wr_addr_s103 : std_logic_vector(9 downto 0);
signal rd_addr_s104 : std_logic_vector(9 downto 0);
signal row_s105 : std_logic_vector(4 downto 0);
signal wren_s106 : std_logic_vector(0 downto 0);


signal ready_s13 : std_logic;
signal done_s14 : std_logic;
signal start_s15 : std_logic;
signal ack_s16 : std_logic;
signal load_done_s17 : std_logic;
signal din_s18 : std_logic_vector(79 downto 0);
signal dout_s19 : std_logic_vector(79 downto 0);
signal addr_s20 : std_logic_vector(9 downto 0);
signal out_addr_s21 : std_logic_vector(7 downto 0);
signal row_s22 : std_logic_vector(3 downto 0);
signal wren_s23 : std_logic_vector(9 downto 0);


signal ready_s108 : std_logic;
signal done_s109 : std_logic;
signal start_s110 : std_logic;
signal din_s111 : std_logic_vector(79 downto 0);
signal dout_s112 : std_logic_vector(79 downto 0);
signal wr_addr_s113 : std_logic_vector(9 downto 0);
signal rd_addr_s114 : std_logic_vector(9 downto 0);
signal row_s115 : std_logic_vector(4 downto 0);
signal wren_s116 : std_logic_vector(9 downto 0);


signal ready_s25 : std_logic;
signal done_s26 : std_logic;
signal start_s27 : std_logic;
signal ack_s28 : std_logic;
signal load_done_s29 : std_logic;
signal din_s30 : std_logic_vector(79 downto 0);
signal dout_s31 : std_logic_vector(79 downto 0);
signal addr_s32 : std_logic_vector(8 downto 0);
signal out_addr_s33 : std_logic_vector(7 downto 0);
signal row_s34 : std_logic_vector(3 downto 0);
signal wren_s35 : std_logic_vector(9 downto 0);


signal ready_s118 : std_logic;
signal done_s119 : std_logic;
signal start_s120 : std_logic;
signal din_s121 : std_logic_vector(79 downto 0);
signal dout_s122 : std_logic_vector(79 downto 0);
signal wr_addr_s123 : std_logic_vector(7 downto 0);
signal rd_addr_s124 : std_logic_vector(8 downto 0);
signal row_s125 : std_logic_vector(3 downto 0);
signal wren_s126 : std_logic_vector(9 downto 0);


signal ready_s37 : std_logic;
signal done_s38 : std_logic;
signal start_s39 : std_logic;
signal ack_s40 : std_logic;
signal load_done_s41 : std_logic;
signal din_s42 : std_logic_vector(79 downto 0);
signal dout_s43 : std_logic_vector(79 downto 0);
signal addr_s44 : std_logic_vector(7 downto 0);
signal out_addr_s45 : std_logic_vector(5 downto 0);
signal row_s46 : std_logic_vector(2 downto 0);
signal wren_s47 : std_logic_vector(9 downto 0);


signal ready_s128 : std_logic;
signal done_s129 : std_logic;
signal start_s130 : std_logic;
signal din_s131 : std_logic_vector(79 downto 0);
signal dout_s132 : std_logic_vector(79 downto 0);
signal wr_addr_s133 : std_logic_vector(7 downto 0);
signal rd_addr_s134 : std_logic_vector(7 downto 0);
signal row_s135 : std_logic_vector(3 downto 0);
signal wren_s136 : std_logic_vector(9 downto 0);



signal ready_s49 : std_logic;
signal done_s50 : std_logic;
signal start_s51 : std_logic;
signal ack_s52 : std_logic;
signal in_a_s53 : std_logic_vector(629 downto 0);
signal out_a_s54 : std_logic_vector(439 downto 0);
signal out_offset_s55 : unsigned(5 downto 0);
signal simd_offset_s56 : std_logic_vector(2 downto 0);
signal op_argument_s57 : sfixed(12 downto -15);
signal op_result_s58 : sfixed(2 downto -8);
signal op_send_s59 : std_logic;
signal op_receive_s60 : std_logic;


signal ready_s139 : std_logic;
signal done_s140 : std_logic;
signal start_s141 : std_logic;
signal ack_s142 : std_logic;
signal din_s143 : std_logic_vector(79 downto 0);
signal dout_s144 : std_logic_vector(629 downto 0);
signal wr_addr_s145 : std_logic_vector(5 downto 0);
signal rd_addr_s146 : std_logic_vector(2 downto 0);
signal wren_in_s147 : std_logic_vector(9 downto 0);

signal input_s62 : sfixed(12 downto -15);
signal offset_s63 : unsigned(5 downto 0);
signal output_s64 : sfixed(13 downto -15);
signal op_send_s65 : std_logic;
signal op_receive_s66 : std_logic;

signal input_s68 : sfixed(13 downto -15);
signal output_s69 : sfixed(13 downto -15);
signal op_send_s70 : std_logic;
signal op_receive_s71 : std_logic;



signal ready_s73 : std_logic;
signal done_s74 : std_logic;
signal start_s75 : std_logic;
signal ack_s76 : std_logic;
signal in_a_s77 : std_logic_vector(439 downto 0);
signal out_a_s78 : std_logic_vector(119 downto 0);
signal out_offset_s79 : unsigned(3 downto 0);
signal simd_offset_s80 : std_logic_vector(0 downto 0);
signal op_argument_s81 : sfixed(12 downto -14);
signal op_result_s82 : sfixed(3 downto -8);
signal op_send_s83 : std_logic;
signal op_receive_s84 : std_logic;



signal ready_s150 : std_logic;
signal done_s151 : std_logic;
signal start_s152 : std_logic;
signal ack_s153 : std_logic;
signal previous_a_s154 : std_logic_vector(439 downto 0);
signal next_a_s155 : std_logic_vector(439 downto 0);

signal input_s86 : sfixed(12 downto -14);
signal offset_s87 : unsigned(3 downto 0);
signal output_s88 : sfixed(13 downto -14);
signal op_send_s89 : std_logic;
signal op_receive_s90 : std_logic;


signal input_s92 : sfixed(13 downto -14);
signal output_s93 : sfixed(3 downto -8);
signal op_send_s94 : std_logic;
signal op_receive_s95 : std_logic;




begin

conv_layer_mc_u0 : conv_layer_mc generic map(
    stride => 1,
    filter_size => 3,
    filter_nb => 10,
    input_size => 30,
    channels => 1,
    dsp_alloc => 1,
    weight_file => "convtest_w0.txt",
    bias_file => "convtest_b0.txt",
    input_int_part => 1,
    input_frac_part => 8,
    weight_int_part => 1,
    weight_frac_part => 8,
    bias_int_part => 1,
    bias_frac_part => 8,
    out_int_part => 0,
    out_frac_part => 8
) port map(
    clk => clk,
    ready => ready_s1,
    done => done_s2,
    start => start_s3,
    ack => ack_s4,
    load_done => load_done_s5,
    din => din_s6,
    dout => dout_s7,
    addr => addr_s8,
    out_addr => out_addr_s9,
    row => row_s10,
    wren => wren_s11
);
bram_pad_interlayer_u97 : bram_pad_interlayer generic map(
    init_file => "~/felix/Git/keragen/convtest_gen/imagedata_7.txt",
    channels => 1,
    channel_width => 9,
    zero_padding => 1,
    layer_size => 28
) port map(
    clk => clk,
    ready => ready_s98,
    done => done_s99,
    start => start_s100,
    din => din_s101,
    dout => dout_s102,
    wr_addr => wr_addr_s103,
    rd_addr => rd_addr_s104,
    row => row_s105,
    wren => wren_s106
);
maxpool_layer_mc_u12 : maxpool_layer_mc generic map(
    pool_size => 2,
    stride => 2,
    input_size => 28,
    channels => 10
) port map(
    clk => clk,
    ready => ready_s13,
    done => done_s14,
    start => start_s15,
    ack => ack_s16,
    load_done => load_done_s17,
    din => din_s18,
    dout => dout_s19,
    addr => addr_s20,
    out_addr => out_addr_s21,
    row => row_s22,
    wren => wren_s23
);
bram_pad_interlayer_u107 : bram_pad_interlayer generic map(
    init_file => "",
    channels => 10,
    channel_width => 8,
    zero_padding => 0,
    layer_size => 28
) port map(
    clk => clk,
    ready => ready_s108,
    done => done_s109,
    start => start_s110,
    din => din_s111,
    dout => dout_s112,
    wr_addr => wr_addr_s113,
    rd_addr => rd_addr_s114,
    row => row_s115,
    wren => wren_s116
);
conv_layer_mc_u24 : conv_layer_mc generic map(
    stride => 1,
    filter_size => 5,
    filter_nb => 10,
    input_size => 18,
    channels => 10,
    dsp_alloc => 1,
    weight_file => "convtest_w1.txt",
    bias_file => "convtest_b1.txt",
    input_int_part => 0,
    input_frac_part => 8,
    weight_int_part => 1,
    weight_frac_part => 8,
    bias_int_part => 1,
    bias_frac_part => 8,
    out_int_part => 0,
    out_frac_part => 8
) port map(
    clk => clk,
    ready => ready_s25,
    done => done_s26,
    start => start_s27,
    ack => ack_s28,
    load_done => load_done_s29,
    din => din_s30,
    dout => dout_s31,
    addr => addr_s32,
    out_addr => out_addr_s33,
    row => row_s34,
    wren => wren_s35
);
bram_pad_interlayer_u117 : bram_pad_interlayer generic map(
    init_file => "",
    channels => 10,
    channel_width => 8,
    zero_padding => 2,
    layer_size => 14
) port map(
    clk => clk,
    ready => ready_s118,
    done => done_s119,
    start => start_s120,
    din => din_s121,
    dout => dout_s122,
    wr_addr => wr_addr_s123,
    rd_addr => rd_addr_s124,
    row => row_s125,
    wren => wren_s126
);
maxpool_layer_mc_u36 : maxpool_layer_mc generic map(
    pool_size => 2,
    stride => 2,
    input_size => 14,
    channels => 10
) port map(
    clk => clk,
    ready => ready_s37,
    done => done_s38,
    start => start_s39,
    ack => ack_s40,
    load_done => load_done_s41,
    din => din_s42,
    dout => dout_s43,
    addr => addr_s44,
    out_addr => out_addr_s45,
    row => row_s46,
    wren => wren_s47
);
bram_pad_interlayer_u127 : bram_pad_interlayer generic map(
    init_file => "",
    channels => 10,
    channel_width => 8,
    zero_padding => 0,
    layer_size => 14
) port map(
    clk => clk,
    ready => ready_s128,
    done => done_s129,
    start => start_s130,
    din => din_s131,
    dout => dout_s132,
    wr_addr => wr_addr_s133,
    rd_addr => rd_addr_s134,
    row => row_s135,
    wren => wren_s136
);
fc_layer_u48 : fc_layer generic map(
    input_width => 490,
    output_width => 40,
    simd_width => 70,
    input_spec => fixed_spec(fixed_spec'(int => 1, frac => 8)),
    weight_spec => fixed_spec(fixed_spec'(int => 1, frac => 7)),
    op_arg_spec => fixed_spec(fixed_spec'(int => 13, frac => 15)),
    output_spec => fixed_spec(fixed_spec'(int => 3, frac => 8)),
    n_weights => 19600,
    pick_from_ram => true,
    weights_filename => "whatever",
    weight_values => reals(reals'( 0.2149530, 0.0095389, 0.1111166, 0.1233901, 0.1717266, -0.0969969, 0.0552405, 0.0860384, 0.1387925, 0.0595221, 0.1157987, 0.0882257, 0.0327046, 0.1285498, 0.1280521, 0.0192293, 0.1140901, 0.0162256, 0.0352322, 0.0403484, 0.0303405, 0.0026690, -0.0068742, 0.0111704, 0.0161444, 0.1559964, 0.1251138, 0.0758125, 0.0981703, -0.0671279, 0.0561959, -0.0586092, 0.0414969, 0.1310353, 0.2299080, 0.0450801, 0.1292331, 0.1526483, 0.0165462, 0.0468746, 0.0349722, -0.1010901, -0.0423811, -0.0796459, 0.1838002, -0.0528305, 0.0142324, -0.0306021, 0.1417059, 0.0447618, 0.1078507, 0.0545914, -0.0401500, 0.1036260, 0.0086952, 0.0088889, 0.0062390, -0.1037199, -0.0600047, 0.0626809, -0.0289324, 0.0610875, 0.0781013, 0.0226872, 0.0146176, -0.0226056, -0.0375533, 0.0324016, -0.0389548, 0.0228771, 0.0898017, -0.0184007, -0.0280840, 0.0131020, 0.0010094, -0.0050012, -0.0498171, 0.0554264, -0.0635130, -0.0586071, 0.1105984, 0.1165285, -0.1980723, -0.0507459, 0.1037367, 0.0730255, 0.1553048, 0.2551782, -0.1054947, 0.0704901, 0.0109695, 0.1969578, 0.2250797, 0.2565585, 0.0817626, -0.1844021, -0.0351138, -0.0158906, 0.2165869, -0.0285433, 0.0332765, -0.2057894, -0.1884436, 0.2026132, 0.1448215, 0.0191223, 0.1387680, 0.2385387, 0.1312052, 0.0425652, -0.0564667, 0.2044180, -0.2105977, -0.0114865, 0.3503435, -0.2756082, 0.0011467, 0.0575665, 0.0064943, 0.0920854, 0.0569069, 0.1488840, -0.0592779, -0.0884504, 0.0862041, 0.0648416, 0.1669873, 0.2213531, -0.0020916, 0.1369014, 0.0458271, 0.2347782, 0.1506993, 0.2433823, 0.1422484, -0.0940610, -0.1723546, 0.0793912, 0.2598021, 0.0753144, 0.0654672, -0.1374128, -0.1040594, 0.0922333, 0.1243162, 0.0421676, 0.1871651, 0.1772649, 0.0891324, 0.0687265, -0.0611514, 0.2081322, -0.1621189, 0.0374418, 0.2749138, -0.2115101, 0.0234102, -0.0872126, -0.0355032, 0.1084775, -0.0146929, 0.0992750, 0.0362255, 0.0298508, 0.1417085, 0.0545119, -0.0186649, -0.0309585, 0.0472688, 0.0794909, 0.0189627, 0.0209592, 0.0584827, -0.0859926, 0.1734718, 0.2214152, -0.0262831, 0.1539500, 0.0342352, 0.0281622, 0.0978196, 0.0641302, 0.1149300, 0.0964129, 0.0761973, 0.1065830, 0.0569699, 0.0370232, 0.0638267, 0.1555289, 0.1428783, 0.0937912, 0.0990565, 0.0594532, 0.0944720, 0.2307579, -0.0771629, 0.0880791, 0.2174948, 0.0215579, 0.0673331, 0.0597854, -0.0463315, 0.1942503, -0.0270705, -0.0281139, 0.2342120, -0.1232101, -0.1320479, 0.2290401, 0.0245070, -0.1093983, -0.0775750, -0.1134888, 0.0837370, -0.0038495, -0.0426198, 0.2411508, -0.0078696, 0.2133640, 0.0575115, -0.0755958, 0.1402902, 0.4384676, 0.1421071, 0.0570157, 0.2268178, -0.0312675, 0.1443339, 0.3990457, 0.0370480, -0.1266562, 0.0543879, 0.2069674, 0.1828734, 0.2002024, -0.0871424, 0.2315755, 0.2161222, 0.0746796, 0.1807910, -0.0486995, -0.0576861, 0.0679277, 0.1294139, -0.0859635, 0.2134576, 0.0000832, -0.0317397, 0.0536612, 0.0172196, -0.0186669, 0.0629640, -0.0783681, 0.0837239, -0.0469428, 0.0817719, 0.0457441, 0.0531505, 0.0437417, -0.0266260, -0.0459630, 0.0909628, 0.0481629, 0.0258416, 0.0118536, 0.0638352, -0.0077420, -0.0417694, -0.0024312, 0.1830197, -0.0836790, -0.0060943, 0.0856343, 0.1934074, 0.0580124, 0.0132292, 0.1366857, 0.0361942, 0.1060068, 0.1307049, 0.0012862, 0.2042811, 0.0838178, 0.1225378, -0.1186724, 0.0505682, -0.0837001, 0.2216204, 0.0943728, 0.1057350, -0.0230773, -0.1281829, -0.0511449, 0.2132953, 0.0160606, 0.2673448, 0.0914931, -0.0287723, 0.1283414, 0.0156265, 0.2371857, 0.2415791, 0.0001850, -0.0129385, -0.1703922, 0.0724498, -0.0625972, 0.0400581, 0.1029179, 0.0939139, -0.1467837, -0.0186173, 0.2536297, 0.1502515, 0.1977101, 0.1857590, 0.0930931, 0.0083272, -0.0076686, 0.1979353, -0.1055420, 0.0684561, 0.0769549, 0.1260012, -0.1480678, 0.0227916, -0.1195581, 0.1644472, 0.1940405, 0.0563370, 0.0268150, -0.0358507, -0.0882061, 0.1287096, -0.0455899, 0.0664386, 0.1330847, -0.0468756, 0.1424174, 0.1069079, -0.0710687, 0.1119290, 0.0031235, -0.1257215, 0.0313911, 0.0716895, 0.0460947, 0.0479687, 0.1374186, 0.0663511, -0.1838419, 0.0958532, 0.0889599, 0.1137180, 0.1799353, 0.1402632, 0.1880081, 0.2133798, 0.0235270, 0.0325615, 0.0570438, -0.0993203, -0.0846650, -0.0788951, -0.0848137, 0.1476005, 0.0062279, -0.1272552, 0.1003162, -0.0258004, 0.0868432, -0.0975145, 0.0768175, 0.0666180, -0.0298739, -0.0372355, 0.0597822, -0.0384823, 0.0088606, -0.0782487, 0.0993932, 0.1432378, -0.0023957, 0.1219289, -0.0080438, 0.0997254, 0.0237937, -0.1163530, 0.1026197, -0.0585502, 0.1008274, 0.2062851, -0.0148296, 0.0345477, 0.0613504, -0.0977356, 0.1213748, 0.0494952, 0.1477299, 0.1378275, 0.1292100, 0.1289798, 0.1912101, 0.1129618, -0.1865616, 0.3030021, 0.1916612, 0.0629863, 0.1299747, -0.0047217, 0.2090874, 0.2281617, 0.1645433, 0.1146196, 0.0178100, 0.0337386, 0.1229954, 0.0931657, 0.0815085, 0.0343134, 0.0806662, 0.0421122, 0.3209148, 0.1633160, 0.0479133, 0.2971745, 0.0926653, 0.0673723, 0.1391150, -0.0729783, 0.0337902, -0.0149062, 0.1499044, 0.1794042, 0.0477222, 0.1219520, 0.1430413, -0.0288464, 0.0927387, 0.1809729, -0.0971993, 0.0232720, 0.3988352, 0.1567653, -0.0505476, -0.0261260, 0.0610141, 0.2111115, 0.0135973, 0.1475370, 0.2154185, -0.0216913, 0.2378640, 0.2130352, 0.0318924, 0.1079730, -0.2173680, 0.2515140, -0.0867896, 0.1462270, -0.0711064, 0.0153622, 0.2058687, 0.2387803, -0.0459229, -0.0388810, -0.1428310, 0.1705836, 0.1185587, -0.0165721, -0.0059123, -0.1832932, 0.3816199, 0.4008062, -0.2616956, 0.3905182, 0.4720702, -0.1690707, -0.0876263, 0.0710234, 0.1947289, -0.2047453, 0.0182906, 0.1307105, -0.0243057, 0.1678538, 0.1354927, 0.0551359, 0.0059859, -0.0577488, 0.2794370, 0.1393692, 0.3540212, 0.0320996, -0.3522376, -0.0697983, -0.0537140, 0.1752933, -0.1481958, -0.0528159, -0.1753761, -0.1335415, 0.0566967, 0.1689524, 0.0402667, 0.1229986, 0.0541515, 0.0664722, -0.1042210, -0.1226066, 0.1758289, -0.1526652, -0.0445802, 0.3777672, -0.3885951, 0.2902862, 0.1338512, -0.0969716, 0.0232866, 0.0767389, 0.0312866, -0.0030267, -0.2145946, 0.0972162, -0.0351145, 0.0304715, 0.0944876, -0.0500789, 0.1034741, 0.0380774, 0.2597741, -0.0147518, 0.1409854, 0.0963850, -0.0549636, -0.0693070, -0.0549658, 0.0533492, 0.0123643, 0.0374218, -0.0818411, -0.0151648, -0.0165146, 0.0321928, 0.0952892, 0.1934236, 0.0254424, 0.0885776, -0.2165439, -0.0281794, 0.0394723, -0.0429591, -0.1900251, 0.1285967, -0.0813443, 0.0842795, -0.2158628, -0.0326722, 0.1378897, -0.0509157, 0.1486267, 0.0132864, 0.1325153, 0.0351053, 0.2344045, -0.0627490, -0.0520579, -0.0618233, 0.2910022, 0.1895111, -0.0767893, 0.0436383, -0.1445236, 0.0277214, 0.3042180, 0.1764989, 0.0564893, -0.0441962, 0.4447573, 0.2851909, 0.2944419, 0.3131101, 0.1838967, 0.0714248, -0.0679312, 0.0691573, 0.2439043, -0.0999673, 0.1725326, 0.3519700, -0.0938588, 0.3922448, 0.2846869, -0.0478876, 0.3231331, -0.2574304, -0.0735464, 0.2122760, 0.1164988, -0.0190222, -0.0340782, -0.0112987, 0.0343971, 0.0225519, 0.1027589, -0.0074442, -0.1756147, -0.1197792, 0.0737163, 0.0114131, 0.0211720, -0.1279679, 0.0045528, 0.0131654, 0.0702988, 0.0331627, -0.0723255, -0.0340449, 0.1617605, 0.0280612, -0.0681802, 0.0288640, 0.1980318, -0.0243412, -0.0403646, 0.0851934, -0.0780333, -0.0039555, 0.1334406, 0.1158854, -0.1050120, -0.0336496, 0.0268874, 0.0955826, 0.0587938, -0.1360784, -0.0410363, 0.0608118, -0.0213011, 0.2792837, -0.0870856, 0.1436989, 0.1442218, 0.3467495, -0.2433292, 0.2202604, -0.1962687, 0.0941692, 0.2825833, -0.1459424, -0.1065909, -0.0281413, -0.0534791, 0.0505372, 0.1123293, 0.1191867, 0.2479287, -0.1596218, 0.3184774, 0.0171047, 0.1462208, 0.2406012, 0.3525361, -0.0451984, 0.0845695, 0.2748735, 0.0442969, -0.0052251, 0.1529491, 0.3088523, -0.3599254, 0.0497125, 0.3152100, 0.2623187, 0.2398119, 0.0822896, 0.2830221, 0.1577007, -0.0780179, 0.2474161, 0.0037491, 0.3014170, 0.3783884, 0.1867528, -0.2002915, 0.2258164, 0.0095973, 0.0975771, 0.1006689, 0.1061653, 0.0191868, 0.2562559, 0.0112711, 0.1839978, 0.1382893, 0.1081401, 0.3528963, -0.0245390, 0.2613134, 0.1031018, 0.2845681, 0.1327966, 0.2613087, 0.1373825, 0.1252876, 0.3223551, 0.0821883, 0.1294325, 0.1743439, 0.0810723, -0.1692714, 0.1417348, 0.3092511, 0.2882398, 0.4055600, -0.0169776, 0.3799770, -0.0536942, 0.0519579, 0.1228539, -0.0219847, 0.2855900, 0.1619733, 0.2112514, -0.1586600, -0.0031646, -0.2110776, 0.1180926, 0.0651365, 0.0124535, -0.1726557, -0.0541247, -0.0223207, 0.1796320, 0.0992658, 0.2099504, 0.1208479, -0.1243740, 0.1663470, 0.0471204, 0.3221792, 0.2061147, 0.0005258, -0.0475033, -0.1525391, 0.1298885, -0.1155267, -0.1744166, 0.0480518, 0.1211077, -0.2213253, 0.1020883, 0.1810327, 0.1300126, 0.1685003, 0.0782781, 0.1150517, -0.0242110, -0.0385910, -0.0232979, 0.1691579, -0.0834911, 0.0087400, -0.0300772, -0.0022185, 0.4428546, 0.1694429, -0.1015083, 0.2875717, -0.0229513, 0.1698840, 0.0807569, 0.0118506, -0.1225642, -0.0290958, -0.0710134, 0.1840827, 0.1000206, 0.3181672, 0.0422843, 0.0342328, 0.1563750, 0.3178539, 0.2293072, 0.0121765, 0.3761014, 0.0861707, 0.0048668, 0.1072557, -0.0416215, 0.1528414, 0.1518032, 0.0577945, 0.3685652, 0.1020111, -0.0756170, 0.1648394, -0.0114091, 0.2257895, 0.0479281, -0.0019347, -0.1940409, 0.1546528, 0.0531214, -0.1244169, 0.1346571, 0.1262165, -0.0142152, 0.2484029, -0.0853981, 0.1370273, 0.1840684, 0.1380555, 0.0366387, -0.0651481, -0.1922279, 0.1834898, 0.0076433, -0.0269425, 0.0568066, 0.0452518, 0.0124177, 0.3163168, 0.1457507, 0.0788811, 0.1810120, 0.1031199, 0.0963593, 0.2160562, -0.0545553, 0.0074590, 0.0499153, 0.1364252, 0.2826516, -0.1018769, 0.1074471, 0.1147052, 0.0222509, -0.0169166, 0.3447673, -0.1296047, 0.1208460, 0.5209471, 0.1429836, 0.0100727, -0.0179959, -0.0120024, 0.1256217, -0.0548513, 0.2093929, 0.0727829, 0.2679097, 0.1013587, 0.2060111, -0.1099712, 0.0229701, 0.1820703, 0.1224120, -0.3369587, 0.0499459, -0.1474651, 0.1074164, 0.3418867, 0.1270311, 0.1584535, -0.0290188, -0.1939000, 0.2894943, 0.1095837, -0.2569828, -0.0332178, -0.1683387, 0.3199672, 0.2433998, -0.3844979, 0.4614383, 0.4750862, -0.2131677, -0.2622935, 0.0878298, 0.1230203, -0.0253027, 0.0913221, 0.0513600, -0.0036774, 0.1247185, 0.0526347, 0.1450718, 0.0766976, 0.0631681, 0.2323439, 0.1418142, 0.2583411, 0.1199625, -0.0737433, -0.0125622, -0.0151468, 0.0998278, -0.0135007, 0.0934319, -0.0036679, -0.0295386, 0.1629389, 0.1455956, 0.1277801, 0.2033244, 0.0279674, 0.1199492, 0.0799451, -0.0307635, 0.1084534, -0.0346897, 0.0326395, 0.1313944, -0.1063633, 0.1651888, 0.1237057, -0.0518178, -0.1037825, -0.0480588, -0.0371308, 0.0764532, -0.2641747, 0.0471103, 0.0837911, -0.0894676, -0.0285011, 0.0663473, 0.1419854, 0.0032698, 0.0247472, -0.0063313, -0.0234962, 0.0459326, 0.0191207, 0.0583974, -0.0744926, -0.0442367, 0.1691439, 0.1777369, 0.0428280, 0.0670938, -0.1407755, -0.1129157, -0.0475103, 0.0651077, 0.0394749, -0.0594980, -0.0859504, 0.0861977, -0.0673771, 0.0848855, -0.0602514, -0.0403327, 0.0541714, -0.1507226, -0.3386909, 0.0625435, 0.0289709, -0.0148374, 0.1573134, 0.2212313, 0.0770504, 0.0374344, 0.2103658, 0.1467035, -0.0414227, 0.0233206, 0.2547907, 0.2307470, -0.0496847, -0.0491510, -0.0882461, 0.0940940, 0.3211919, 0.3203582, 0.1655684, 0.1417488, 0.3685315, 0.0697410, 0.0682896, 0.2923319, 0.1056199, 0.1084238, -0.0188472, 0.2402674, 0.2522778, -0.1775371, 0.2694940, 0.3148413, -0.0169354, 0.3145969, 0.3121287, 0.0099629, 0.2331669, -0.2623610, -0.0383441, 0.3721249, 0.2901430, -0.0241519, -0.0850862, -0.0188259, -0.1683051, 0.0146718, -0.0210358, -0.0488917, -0.1975433, -0.0566260, 0.0356904, -0.0081287, -0.0396791, -0.0904655, 0.0266475, -0.0129790, 0.0372019, -0.0023098, -0.1635157, 0.0340111, 0.0541915, 0.0229540, 0.0252658, -0.0233519, -0.0516774, 0.0197546, -0.0567444, 0.0517851, -0.1102361, -0.1017384, -0.0007396, 0.0444043, -0.0955964, -0.0142142, -0.0570459, -0.0084899, -0.0314724, -0.1659573, -0.1641852, -0.0155801, 0.0273699, 0.2453142, -0.0996215, 0.3686859, 0.1512076, 0.3570903, -0.2699683, 0.0983864, -0.2704393, 0.1185642, 0.1056216, -0.2662651, 0.0002002, -0.0613222, 0.0180280, 0.3125870, 0.1202066, 0.4105566, 0.0058855, -0.0792259, 0.3728981, -0.0052109, 0.0813550, 0.3856576, 0.0647099, -0.1437241, -0.0286059, 0.2235649, -0.1037925, -0.2910367, -0.0978450, 0.1896767, -0.2480109, -0.0391958, 0.2193068, 0.4572823, 0.1767853, 0.1598027, 0.1538137, 0.1126339, -0.0305019, 0.0925514, 0.0139894, 0.2350146, 0.2519253, 0.1634486, -0.3512279, 0.2577907, -0.2106382, -0.0154551, 0.2113916, -0.2082684, -0.1431016, 0.1271403, -0.0600886, 0.0051178, 0.0275758, 0.1687271, 0.3377366, -0.1989341, 0.2890068, 0.0455297, 0.2201870, 0.1828212, 0.3572214, -0.1073718, -0.0316827, 0.3194328, 0.2168420, -0.1451489, 0.0887082, 0.1321670, -0.4356401, 0.0042125, 0.2682260, 0.4420550, 0.2782223, -0.0262157, 0.2362454, 0.1059305, 0.0534367, 0.1643357, -0.1557386, 0.0905718, 0.1135802, 0.1813710, -0.1232724, -0.0332152, -0.0249622, 0.0884536, 0.0548620, -0.0804684, -0.1521379, -0.1228062, 0.0820028, 0.1426936, 0.1264658, 0.1684360, 0.0030709, -0.1642561, 0.1861431, 0.0479751, 0.0771139, 0.1296835, -0.0095927, 0.0244704, -0.0783176, 0.0436687, -0.0771413, -0.0541669, 0.0830828, 0.1294769, -0.1959650, 0.0267873, 0.1970079, 0.0623626, 0.0010024, -0.0163933, 0.0623969, -0.0577607, 0.0340275, -0.0425202, 0.1116248, -0.1138099, -0.2033928, 0.0761621, -0.1538746, 0.3771547, 0.2166148, -0.0142368, 0.4306993, -0.1664831, 0.2925543, 0.2583723, 0.3694691, -0.1332999, -0.0247300, -0.0733257, 0.0818254, 0.1095550, 0.3010369, 0.0028603, 0.0955295, -0.0263316, 0.1656586, 0.1805131, 0.0777908, 0.5633604, 0.2905794, -0.1933962, -0.1420352, 0.0094614, 0.0832415, 0.0346121, -0.1383419, 0.2520709, 0.0130659, -0.1000184, -0.2229570, 0.1143126, 0.1849978, -0.0912579, -0.0457193, -0.2036412, 0.0123901, -0.0430234, 0.1314235, 0.1459944, 0.0773276, -0.1101249, 0.1451781, -0.0284119, 0.1089119, 0.0080570, 0.1509086, -0.0142149, -0.0072540, -0.1468788, 0.1336221, 0.1444654, -0.0751171, 0.0616084, 0.0055866, 0.0247437, 0.1808167, 0.1725744, 0.0544102, 0.1602872, -0.1250546, 0.0812312, 0.2688326, -0.0593711, 0.0632001, 0.1260230, 0.0447072, 0.2124584, 0.0472823, 0.0362826, 0.0036756, 0.0017072, -0.0214394, 0.2203430, 0.1182514, -0.0907249, 0.3654732, 0.0659658, 0.0377349, 0.0605109, 0.2062401, 0.1027366, -0.1316564, 0.2215926, 0.0183718, 0.2888494, 0.1633128, 0.2219604, 0.0267131, -0.1167876, 0.1636900, 0.1001497, -0.4532818, 0.0573699, -0.1458062, -0.0074003, 0.3177846, 0.3278655, 0.1997668, -0.0310655, -0.0239760, 0.2883094, 0.2034065, -0.2377174, 0.0427627, -0.1282319, 0.3689675, 0.1597106, -0.4135949, 0.2568038, 0.3877467, -0.1077470, -0.2969342, 0.0991749, 0.0768272, -0.0949462, 0.0977010, 0.0600177, 0.0681945, 0.0257871, 0.1776248, 0.0046607, 0.0552799, 0.1174122, -0.0546125, 0.0828725, 0.0200829, 0.1137619, 0.0384712, -0.0433366, 0.1093666, 0.0105579, -0.1406625, 0.0278762, 0.0060948, -0.0472769, 0.1586293, 0.1232023, 0.1473748, 0.0069857, 0.0066044, 0.1809992, 0.1711858, -0.0124215, 0.0199426, 0.0579956, 0.1721898, 0.0234651, -0.1025922, 0.0609861, 0.1527800, 0.0302290, -0.1188576, 0.0829669, -0.0029432, 0.0281144, -0.2313237, 0.0988757, 0.0183805, -0.0144775, -0.0517358, 0.0356748, 0.1194081, 0.0291776, 0.0418323, -0.0603749, 0.0084034, 0.0051887, 0.0569994, 0.0518861, -0.0295774, -0.0135580, 0.0745530, 0.1027738, 0.0619366, 0.0450006, -0.1079522, -0.0933899, 0.0294397, 0.0417527, 0.0944061, -0.0280485, 0.0336423, 0.0367513, -0.0288882, 0.0530368, -0.0366569, -0.1041351, 0.0532712, -0.1498996, -0.3093068, 0.0469533, 0.0320854, 0.0963431, 0.1444975, 0.0559587, -0.1287671, 0.0922104, -0.0606052, 0.2710409, 0.2017123, 0.2071430, 0.0630390, -0.0908800, 0.0637866, 0.1731404, 0.1459684, 0.1557021, 0.0502490, 0.0305933, 0.1565381, 0.2290854, 0.1180066, -0.1521063, -0.1239742, 0.0504445, -0.1637312, 0.0542071, 0.0367313, 0.1093922, 0.2692720, -0.2237026, -0.2495023, 0.0349297, 0.2045231, -0.0462858, -0.0816661, -0.0081951, 0.0312860, 0.0642389, -0.1532175, 0.1521617, 0.1460089, -0.0178795, -0.0692209, 0.0062144, -0.0607681, -0.0157347, -0.0166183, -0.0518000, -0.1470823, -0.0439233, -0.0100981, -0.0024908, -0.0652318, -0.1271240, -0.0070322, -0.0256049, 0.0307142, 0.0083702, -0.0332041, -0.0666506, 0.0328286, -0.0043935, 0.0550052, -0.0008152, -0.1087980, -0.0865793, -0.0487966, -0.0199873, -0.0468246, -0.0604844, -0.0210145, 0.0120836, -0.1007641, 0.0130124, -0.0615981, -0.0312450, 0.0280205, -0.0903696, -0.1145770, -0.0019263, 0.0022143, 0.4850509, 0.0217302, 0.3967576, 0.3492154, 0.3530502, -0.1570234, -0.0713632, -0.1413493, 0.1648858, -0.1217419, 0.0902551, 0.0513022, 0.1276352, 0.0403671, 0.3201049, 0.0761786, 0.3781380, -0.0524102, -0.0192527, 0.0594625, -0.0607390, -0.0615131, 0.1331367, 0.1007782, -0.0119037, 0.0602376, -0.0859305, 0.1386817, 0.0184476, -0.1262499, 0.0966481, -0.0955113, -0.1554986, 0.3961294, 0.2960218, -0.2111461, 0.1813444, 0.4071540, -0.1451227, -0.1283475, 0.2163427, -0.0946637, 0.3803751, 0.3106565, 0.2893083, -0.3657541, 0.1342276, -0.2236611, 0.1459258, 0.0753820, -0.1657415, -0.0415240, -0.0290612, -0.0048295, 0.1019979, 0.0082891, 0.3882743, 0.1720542, -0.1315293, 0.1050340, -0.0261672, 0.1131398, 0.1724611, 0.0292712, -0.0569809, -0.0438668, 0.1750905, 0.0402557, -0.1218450, -0.0773178, -0.0025926, -0.2734712, -0.0380548, 0.2729954, 0.3220600, 0.1538679, 0.1499946, 0.2723689, -0.1846121, 0.0475688, 0.2652417, 0.0254267, 0.2085707, 0.1464478, 0.2121006, -0.0686728, -0.0949178, -0.1553867, 0.0871544, -0.0236351, -0.1724905, -0.2906582, -0.0533344, -0.2257981, 0.2837715, 0.0874950, 0.2790709, 0.0792354, -0.0825000, 0.2816361, -0.0779002, 0.0172877, 0.2704493, -0.0271767, -0.1262479, -0.1029293, -0.0052950, 0.1151780, -0.1329857, -0.0686005, 0.1685027, -0.3037978, 0.0566177, 0.2504008, 0.1590370, 0.0650786, -0.0282849, 0.1345307, 0.0478902, 0.0199975, 0.1184906, 0.1303681, 0.0527915, -0.3805373, 0.0268084, -0.1553077, 0.3767080, 0.2794770, 0.1119720, 0.4414468, -0.0857842, 0.2263048, 0.1483803, 0.1248535, 0.0853349, 0.0709441, 0.0248145, 0.1975419, 0.0153603, 0.3530556, -0.0037897, -0.0677673, 0.0517736, -0.0425523, -0.1562720, 0.2427272, 0.3706900, 0.3576551, 0.0012694, -0.1601628, 0.0945347, 0.0775575, 0.0325806, -0.3267059, 0.0634403, 0.1773144, -0.2944409, -0.3326941, 0.1682915, 0.2587627, -0.1158790, 0.0133297, -0.0303780, -0.1043573, -0.0760406, 0.1846867, -0.1164768, -0.0696744, -0.1645144, 0.2397615, -0.0035899, 0.0013989, -0.1393032, -0.0967053, 0.1061809, 0.1175702, 0.0330038, -0.1217443, -0.0156526, 0.3253031, 0.1117772, 0.1293079, 0.2777102, -0.0148640, 0.0772717, -0.2038246, 0.0384687, -0.0238880, -0.0518577, 0.1286583, 0.1583682, -0.1071370, 0.2218993, 0.0418893, 0.0438211, 0.1913688, -0.2144155, -0.1152171, 0.1003521, 0.1361077, 0.1828170, 0.1400884, -0.0359603, 0.3178477, 0.0448109, 0.1106839, 0.0635125, 0.1115829, 0.1234340, -0.1366198, 0.2649170, 0.0110936, 0.2331177, 0.1332410, 0.1881103, 0.0848447, 0.0062509, 0.1508083, 0.1519573, -0.5386562, 0.0820916, -0.0586640, -0.0630052, 0.3147960, 0.3768571, 0.0969124, -0.0289366, 0.0144129, 0.2058968, 0.2712053, -0.2595915, 0.1263113, -0.0455172, 0.3832319, 0.1438449, -0.4013936, 0.1630900, 0.3029585, -0.2238951, -0.4043575, 0.0852257, 0.0432288, -0.1548639, 0.0743772, -0.0066570, 0.1130733, 0.0209547, 0.0886149, -0.0360947, 0.0316638, 0.1455290, -0.0569648, 0.0935530, 0.0874417, 0.1393027, 0.0723075, -0.1041646, 0.0479526, 0.0280954, -0.1390102, 0.1266385, -0.0536627, -0.0195961, 0.1318153, 0.2278032, 0.0760013, 0.0316679, 0.0229225, 0.1582822, 0.2555178, 0.0006391, 0.0875751, 0.0420167, 0.1596179, -0.0242736, -0.1026909, 0.0836216, 0.0466390, -0.0007900, -0.2841563, 0.0648122, 0.0528776, 0.0163741, -0.1340922, 0.0827121, -0.0678751, 0.0531475, -0.0068101, 0.0664663, -0.0021034, -0.0033029, 0.0607141, -0.0211043, 0.0759059, 0.0230872, 0.0169462, 0.0557711, -0.0294815, -0.0017805, 0.0228971, 0.0240429, 0.0493585, -0.0127147, -0.1325674, 0.0136944, 0.0382249, 0.0904236, 0.1186496, 0.0100452, -0.0865959, -0.0542816, -0.0112025, -0.0270228, -0.0223584, -0.0946329, 0.0131665, -0.0294774, -0.1643861, -0.0364634, -0.0019394, 0.0864647, 0.1357589, 0.3641630, -0.2974188, 0.1529263, 0.2331745, -0.0837017, 0.1199526, 0.1383965, -0.0267045, 0.1495847, 0.1263434, -0.0253058, -0.1978934, 0.1294329, 0.2684766, 0.2263647, 0.2328101, 0.1544055, 0.1806472, 0.1941597, -0.1442459, 0.1866243, -0.1604586, -0.2036225, 0.1271563, -0.2436731, 0.2583429, 0.0579788, -0.3547532, 0.2132286, 0.0706477, 0.0368014, -0.2035739, -0.0994118, 0.2147378, -0.0006563, -0.1847235, 0.3395126, 0.1515856, -0.0984245, -0.0635702, -0.0556464, -0.0327250, 0.0117613, 0.0096193, -0.0894889, -0.1010372, -0.0450259, -0.0415269, 0.0230500, -0.0308264, -0.1335748, 0.0113295, -0.0706666, 0.0071519, 0.0155301, -0.1108538, -0.0577093, -0.0113210, 0.0274213, 0.0435027, -0.0385077, -0.0850912, -0.0149595, -0.0664022, -0.0071713, -0.0755621, -0.0421243, 0.0374948, 0.0110363, -0.0532132, -0.0069134, -0.0246398, -0.0307646, 0.0023659, -0.0901181, -0.0824011, -0.0133441, -0.0237661, 0.3069631, 0.2157989, 0.1193626, 0.2823995, 0.2493380, -0.0312675, 0.0221646, 0.0589716, 0.0041878, -0.1413508, 0.1677275, 0.0404436, 0.3380447, 0.1739465, 0.1898560, 0.2116216, 0.1771614, -0.0222020, 0.1859987, 0.0089609, 0.2050938, -0.0936627, -0.0024961, 0.3062850, 0.2094699, 0.2909583, 0.0090732, 0.2468807, 0.2568920, 0.1768045, 0.0287384, -0.0349046, -0.1482788, 0.3181733, 0.0859459, -0.2307869, 0.0543157, 0.3853920, 0.0181300, -0.3073878, 0.2822037, 0.0888137, 0.3804382, 0.3251941, 0.2542326, -0.3763399, 0.0690496, -0.0846200, 0.1362360, -0.1215139, -0.1329488, 0.0037304, 0.2007703, -0.0311744, 0.1318991, -0.0781032, 0.3380690, 0.2459732, -0.0593530, -0.0633760, -0.0817713, -0.0036118, 0.0857466, 0.2019586, -0.0678388, 0.0370562, 0.0571967, 0.1128844, -0.1213135, -0.1668136, -0.0743733, -0.2450805, -0.1816639, 0.2828136, 0.3209653, -0.0836936, 0.1055748, 0.3344536, -0.1662454, -0.1901221, 0.3915316, 0.1108264, 0.4383993, 0.2571469, 0.3073676, -0.0327123, -0.3428818, -0.0094863, 0.2320128, -0.2814648, -0.0060002, -0.0687005, 0.0828885, -0.0804398, 0.3761606, 0.0661478, 0.4705070, 0.0440380, 0.0336820, -0.3007895, -0.0593819, -0.2655781, 0.1099499, 0.0237353, -0.0183892, -0.0020401, -0.3503944, 0.1740518, 0.0076073, -0.2293779, 0.0143080, -0.0682655, -0.2095584, 0.2404175, 0.0014891, -0.3371521, 0.2684939, 0.3235183, -0.1614012, -0.2524880, 0.1041930, 0.0837077, 0.1056295, -0.0407762, 0.0840839, 0.1086415, -0.0119888, 0.0637271, -0.0756193, 0.1698880, -0.0607590, 0.1105657, -0.0187792, -0.1071192, 0.1024678, 0.1140567, 0.0449316, -0.0011987, 0.0581245, 0.4806489, 0.1954779, -0.0047700, 0.0463234, -0.0094012, -0.1873711, 0.1340233, 0.0098090, 0.2035060, 0.1014874, 0.0261710, 0.2588352, -0.0032336, 0.0694549, -0.0751565, 0.0259344, 0.2711973, -0.1779289, -0.1957234, 0.2881967, 0.2295776, 0.0039971, -0.0808847, 0.0963160, 0.0088663, 0.0417147, 0.1855941, -0.1572899, -0.0996460, 0.0126045, 0.2483573, 0.0299198, -0.1666428, -0.3759750, -0.0563731, 0.1523286, 0.1488666, 0.1384621, -0.0401007, -0.0921895, 0.3014198, 0.0879605, 0.1579864, 0.2967673, -0.0591701, 0.0532666, -0.1800922, -0.0064570, -0.1172958, -0.1607317, 0.2034387, 0.1974815, -0.1543543, 0.2477176, 0.1614583, -0.0539544, 0.0841135, -0.1175130, -0.0033990, 0.0272905, 0.1710488, 0.0526371, 0.0077460, -0.0804619, 0.2891450, -0.0220004, 0.3398809, -0.2842025, 0.0995968, 0.0575201, -0.1515701, 0.4900871, 0.0138380, 0.1895829, 0.1853745, 0.2411745, 0.1522138, -0.0126066, -0.0693756, 0.1389021, -0.3249972, 0.1035826, -0.1440948, -0.0714337, 0.1736089, 0.3518269, -0.1506442, -0.2696497, -0.0145340, 0.3118067, 0.2032199, -0.1663119, 0.2112765, -0.0657971, 0.3024314, 0.0567723, -0.2852938, 0.2881804, 0.3754191, -0.1689179, -0.2390516, -0.0034779, -0.1915483, -0.2056026, 0.1412984, -0.1517210, 0.3540187, -0.1284498, 0.0344797, 0.1812029, -0.0123689, 0.3751964, 0.2493137, -0.0517925, 0.3853112, 0.0447463, 0.0330465, -0.1403798, -0.1244858, 0.3105347, -0.2693536, 0.3074374, 0.1203527, -0.0046938, 0.0423342, 0.3567407, 0.0420978, -0.1589449, -0.2046570, 0.2302341, 0.3552574, -0.1004930, 0.2148826, 0.0279262, 0.3063662, -0.0615290, -0.1365864, 0.2575597, -0.0004030, -0.1138930, -0.1762630, 0.0439315, 0.0805102, 0.0972112, -0.0479263, 0.0949645, -0.0328710, 0.1144061, 0.0346304, 0.1911131, -0.1161640, 0.1390702, 0.0533270, 0.0714240, 0.0998493, -0.0213827, -0.0146670, 0.0907317, 0.0280563, 0.0093542, -0.1504923, 0.0646990, 0.1365716, -0.0505271, -0.1095288, 0.0946900, 0.0688590, 0.1122239, 0.0382925, 0.0262740, -0.1211832, -0.1127225, 0.1064200, -0.0480846, -0.0062540, -0.0472716, -0.0032786, 0.1269087, -0.0258748, -0.1547047, -0.0362981, 0.1342601, 0.1964560, 0.2758135, -0.0638770, 0.2613407, 0.2495826, -0.2118556, 0.0453201, 0.1214711, -0.0075962, 0.1255161, 0.2166172, 0.0822159, -0.1726658, 0.1602024, 0.2197942, 0.3341610, 0.0167436, 0.1506398, 0.1659524, 0.2307834, -0.1015775, 0.0372179, -0.0989062, -0.1333303, 0.0342777, -0.0716029, 0.3377089, 0.2135413, -0.1487232, 0.1810634, 0.1199104, 0.0060103, -0.0387748, -0.0706432, 0.1231009, 0.0328477, 0.0247312, 0.2071536, 0.1025914, 0.0358190, -0.0906066, 0.0055435, -0.0047334, 0.0374955, -0.0187128, -0.0363723, -0.0256329, 0.0320091, -0.0555351, 0.0373535, -0.0374271, -0.0831144, 0.0517255, -0.0083445, -0.0037802, 0.0620042, -0.0448894, -0.0209062, -0.0159334, 0.0001488, 0.0644456, 0.0037892, -0.1133495, 0.0392944, -0.0286853, 0.0151824, -0.0943647, -0.0653796, 0.0264879, -0.0141506, 0.0029775, -0.0174946, 0.0339007, -0.0806482, -0.0237932, -0.0171816, -0.0242062, -0.0621442, -0.0517403, 0.2323872, 0.1419313, -0.1465179, 0.2277790, 0.1669974, -0.0810508, 0.3388599, 0.1017206, -0.0458758, 0.1807791, 0.1685863, 0.2388498, 0.2615982, 0.2559305, 0.0303650, 0.1028583, -0.0388437, 0.2533841, 0.1438879, 0.2511033, 0.1429527, 0.1117165, 0.0164318, 0.3641406, 0.3614189, 0.3319418, 0.3928981, 0.2138954, 0.2685322, 0.4052018, 0.1399229, 0.0287290, 0.1077364, 0.1536800, 0.1147237, 0.1701400, -0.0523410, 0.3218786, 0.1382348, 0.0740785, 0.2392353, 0.0697784, 0.3267950, 0.2180615, 0.2692100, -0.0898943, 0.0710541, 0.0502826, 0.1327636, -0.0687263, -0.0003350, -0.0326145, 0.0771459, 0.0571636, 0.0862131, 0.0460218, 0.2680722, 0.1706961, 0.0822701, -0.0422397, 0.0100900, -0.0824556, 0.0778557, 0.1215133, 0.0590353, 0.0952849, 0.0546436, 0.2090469, 0.0703658, -0.0281739, -0.0681837, -0.0129050, -0.0918507, 0.2650686, 0.1816440, -0.0273577, 0.1218542, 0.2107930, -0.1414040, -0.1465368, 0.4278079, -0.1618496, 0.5607112, 0.4241666, 0.3896280, -0.1916061, -0.0715625, -0.0632519, 0.3985334, -0.2297282, -0.0689049, 0.1500371, 0.0126563, 0.1203818, 0.3377396, -0.0768417, 0.5261419, 0.2490222, 0.0498046, -0.2975757, -0.0461126, -0.0591846, 0.2063152, 0.1411226, 0.0020801, 0.0737753, -0.1694992, -0.1064073, 0.0941711, -0.1859134, -0.2005170, 0.0497585, -0.2059574, 0.5001439, 0.4015422, -0.0981732, 0.3439936, 0.4218141, -0.3307092, -0.2757021, 0.0878917, 0.2397215, 0.1897326, -0.0534993, 0.1112542, 0.2304116, -0.1874570, -0.1266818, -0.0174239, 0.0474664, 0.2350923, -0.0871002, -0.1942417, -0.1391577, 0.1533885, 0.3087844, 0.3245050, -0.0215125, 0.1386388, 0.3481454, 0.1705630, -0.0155601, 0.1700164, -0.0736806, -0.1631857, -0.0762276, -0.0383697, 0.2728873, 0.0347303, 0.0875799, 0.3194328, -0.0169331, 0.0781405, 0.0663091, -0.1403520, 0.1472666, -0.0641559, -0.0167092, 0.1984526, 0.2268820, 0.0390509, -0.1340374, -0.0449268, 0.0104802, 0.1225045, 0.0955162, 0.0046247, -0.0400700, 0.1324999, 0.2364426, 0.0432442, -0.1438576, -0.0685473, 0.0068142, 0.2028538, 0.0849189, 0.1323058, 0.0337462, -0.0236949, 0.1939333, -0.0468676, 0.0325357, 0.1554130, -0.0761589, 0.0973191, -0.0611967, 0.1020082, -0.1241846, -0.0554657, 0.0594733, 0.0875923, -0.0636936, 0.1573743, 0.0551387, -0.0956780, -0.0671570, -0.0435361, 0.0380698, 0.0537970, 0.0448854, -0.0521996, -0.2369584, -0.0405708, 0.2029717, -0.0056329, 0.2853420, -0.0355832, -0.1659716, 0.1294141, -0.0407460, 0.4493916, 0.0760518, 0.0041045, 0.3918752, -0.0410624, 0.0836307, 0.0960474, 0.0084320, 0.0165848, -0.0058712, 0.3673860, 0.0822787, 0.0884236, 0.2010736, 0.2200881, 0.0579907, 0.0512636, -0.2098493, 0.2324380, 0.1973908, -0.0048452, 0.0422814, 0.1434936, 0.3253175, 0.1134416, -0.0827738, 0.1024022, 0.1016257, -0.1369868, -0.1715058, -0.0153915, -0.1145305, -0.0715239, 0.1022407, 0.0053967, 0.0153506, -0.0422208, -0.0175597, 0.0774758, 0.1020648, 0.1396623, -0.0667186, -0.0101504, 0.1065758, 0.0523403, 0.0615823, 0.0759158, -0.0053310, -0.0275992, 0.0553177, 0.1812261, 0.0239260, 0.1372707, -0.0854726, 0.1495729, -0.0050736, 0.1055653, -0.1450118, 0.1368474, 0.1296126, -0.0459409, 0.0211391, 0.0246702, 0.1445398, 0.0008139, 0.0584413, 0.0312588, 0.0473874, -0.2238803, -0.0799818, 0.1599394, -0.0977180, 0.0996267, 0.0046370, 0.2352460, 0.0801618, 0.0227763, 0.0392734, 0.3008272, -0.1887791, 0.4076603, 0.3012338, -0.0041065, 0.5125046, -0.0375986, 0.0130692, 0.2728217, 0.0858064, 0.1469087, -0.3119160, 0.2235474, 0.2756298, -0.0753598, -0.0451052, 0.2307552, 0.1663138, 0.0327420, -0.2260915, 0.1748031, -0.0194945, -0.2146612, 0.2990836, -0.0353264, 0.1548914, -0.0479015, -0.0980975, 0.3911905, 0.1717200, -0.3582246, -0.1425584, 0.1913351, 0.0647970, 0.1248683, -0.0135232, 0.1587137, -0.0327957, 0.0516642, 0.0487478, 0.1300193, 0.0678678, 0.1008819, 0.1127217, 0.1894726, 0.1833096, 0.1685163, 0.0163585, 0.1351958, 0.1519883, 0.0561561, -0.1122700, 0.1988830, -0.0718803, 0.0182720, -0.0420119, 0.1113176, 0.1080725, 0.1424666, -0.0138185, 0.0129871, -0.0816522, -0.0327560, 0.0717611, -0.0523908, 0.0813198, 0.1475136, -0.1070476, 0.1483494, 0.1324593, -0.0737747, 0.0529464, 0.1223975, -0.0586084, 0.0818283, 0.0795073, 0.1154106, 0.0489560, 0.0182135, 0.0567481, 0.1730624, -0.0620499, 0.1198122, -0.0111635, 0.0146219, 0.0962192, 0.0489687, 0.0234836, 0.1089474, 0.0638195, -0.0461251, -0.0996538, 0.0678743, 0.0352167, -0.0115372, -0.0866888, 0.1290049, 0.0533972, 0.0146938, -0.0842977, 0.1399009, 0.0582250, -0.0299533, 0.0724415, 0.0134076, 0.0990595, -0.0714128, -0.0752717, 0.1616056, 0.0799574, -0.1031687, -0.0822036, 0.1828551, 0.0489282, 0.1422513, 0.0598827, 0.1342497, -0.0231456, 0.2448006, 0.1061848, 0.1433685, 0.1076034, 0.0930006, -0.0203820, -0.0149655, 0.0750174, 0.1762311, 0.1048688, 0.1098160, 0.2335350, 0.0177789, 0.1932102, 0.0242030, -0.0405515, 0.0965514, 0.1895275, 0.0800052, 0.1570069, 0.1559977, 0.1224945, 0.2000250, 0.1407050, 0.1276299, 0.0031205, 0.0463696, 0.0858793, 0.0185055, 0.2628644, 0.0941832, 0.0878405, 0.2139909, 0.2149854, 0.1987004, -0.1218234, 0.3719762, 0.2027194, 0.1564568, 0.1087354, -0.0849658, 0.0074017, 0.3096789, -0.0234460, 0.1033068, 0.0343669, -0.0267032, 0.0435195, 0.2735942, 0.0805151, 0.3303627, -0.0074658, 0.1118155, 0.0420100, 0.0497345, -0.0248778, 0.1865222, -0.0128289, -0.0413902, -0.0307698, -0.0480559, 0.0070862, -0.0134856, -0.1360524, 0.0591373, 0.1170994, -0.0950306, 0.3427565, 0.3026779, -0.0553148, 0.2984990, 0.2159012, -0.0682403, -0.1339646, 0.4041953, 0.1219389, 0.4463297, 0.3655259, 0.2433482, 0.0044783, -0.0474428, -0.0274736, 0.1762285, -0.1089574, -0.0609343, 0.1027458, 0.1584288, -0.0187666, 0.2242848, -0.0063618, 0.3562397, -0.0943527, 0.1746697, -0.0705759, -0.0636187, -0.0241727, 0.2732326, 0.0472273, -0.0241945, -0.0357326, -0.0232535, 0.2060141, -0.0099472, -0.0242307, 0.0631177, 0.1134377, -0.1020714, 0.2982357, 0.3193496, -0.1111147, 0.2499433, 0.2348252, -0.1439030, -0.1027882, 0.0510242, 0.0932997, -0.0046569, 0.0682612, 0.0400279, 0.0763014, -0.0213415, 0.1377774, 0.1218921, 0.1879768, -0.0076900, -0.1186121, 0.1307864, -0.0270968, 0.1664265, 0.1636876, 0.1579181, 0.1468006, -0.0725682, 0.2218471, 0.0421020, 0.0244112, 0.1185123, 0.0658224, 0.2044292, -0.0247086, 0.0368701, 0.1858813, -0.1295982, 0.1241023, 0.1958453, -0.0245911, 0.1469570, 0.1210308, -0.0511902, -0.1253027, -0.0027145, 0.0052058, 0.1538877, 0.0665120, 0.0638640, 0.0384785, -0.0640823, -0.0318049, 0.0053636, -0.0378662, -0.0528263, 0.0078323, -0.0813265, 0.0018115, 0.0038527, 0.0513228, 0.1082183, 0.1211587, 0.1518740, 0.0808268, -0.0328890, -0.0591297, 0.1199078, -0.0294258, 0.0012861, -0.0838913, 0.0035796, 0.0748833, 0.1358871, -0.0869272, 0.0513766, 0.0599465, 0.0604732, 0.0482590, 0.0108306, 0.0557847, -0.0659449, 0.0535566, 0.1168774, -0.0582178, 0.1048291, -0.0804566, -0.0289390, -0.0080243, -0.0176704, 0.0904088, 0.0723411, -0.1986012, -0.0460098, 0.0308657, -0.0998080, -0.0318356, -0.0063813, 0.0060154, 0.0856242, 0.0648287, 0.0146840, -0.0968883, 0.1508152, 0.1156606, 0.2070063, -0.1609993, 0.1595534, 0.0544974, 0.0638160, 0.0509230, 0.1672986, -0.1147181, -0.0039447, -0.1142261, -0.0335534, 0.1286641, -0.2078166, -0.1115326, 0.2232435, 0.0697195, 0.0546631, -0.0315463, -0.0121693, -0.0294956, -0.0602348, -0.1840457, -0.0176942, 0.1537512, -0.0841249, 0.2703980, -0.2871484, 0.0888114, -0.1174790, -0.0374545, 0.1543091, 0.2622940, -0.1986819, 0.1458390, 0.0054302, 0.2292681, 0.2093826, 0.5394033, 0.0844931, -0.0029484, -0.1301820, -0.1687539, 0.4213130, 0.1375983, -0.1370055, 0.0022594, 0.0284328, 0.1162877, 0.4550416, -0.1886410, 0.2731154, 0.3120990, -0.1597080, 0.0142541, -0.0947139, 0.1361814, 0.0494362, 0.1638090, 0.2910708, -0.2569810, -0.1567438, -0.0776057, -0.1562835, 0.2967732, -0.1810051, 0.1558775, -0.0719430, -0.0354606, -0.0747732, -0.1396018, 0.0921680, 0.3041607, -0.1542332, 0.2343047, -0.0529473, 0.0875425, 0.0750536, 0.3806210, 0.0349882, -0.0302163, -0.1646972, -0.1631730, 0.2099273, 0.0897051, -0.1019688, -0.0616720, 0.1610890, 0.0834844, 0.3727986, -0.1760506, 0.1597991, 0.2231502, -0.1582156, -0.0303630, 0.0490440, 0.1817803, 0.0470174, 0.0974817, 0.1835119, -0.2993023, -0.0114395, -0.0981258, -0.1387108, 0.3401086, 0.1660604, 0.0843516, -0.1263487, 0.1544285, 0.0676707, 0.1691136, 0.3223242, 0.0372214, -0.1258503, 0.4843851, -0.0625522, 0.0250935, -0.0345976, -0.0949027, -0.0340526, -0.0112218, -0.1950977, 0.1933897, 0.0607739, 0.4528253, 0.1083004, -0.0731770, 0.1190713, 0.3811452, 0.1450671, 0.0150481, 0.2809223, 0.0819638, -0.0353105, 0.4188692, 0.1107902, -0.1281293, 0.1886043, 0.1113319, 0.2948469, 0.3133722, -0.1090638, 0.1191058, 0.1926801, 0.1331724, 0.0380944, 0.1287026, -0.2620308, -0.1109472, 0.0463405, 0.0121197, -0.0353545, 0.0429014, -0.1646242, 0.1761493, -0.1915461, 0.0342740, 0.0258552, 0.0615670, -0.0473496, -0.0012529, -0.1973598, 0.0718360, 0.1405452, 0.1791636, -0.0019171, -0.2223721, -0.0449375, 0.1867590, 0.0369709, -0.0328588, 0.1274591, 0.0176897, 0.0011980, 0.1634228, 0.1164389, -0.1153734, -0.0602833, -0.0898041, 0.1273479, -0.1086954, -0.1349803, -0.0941241, 0.0808337, 0.1105300, 0.1308056, 0.0432280, 0.1601620, 0.1531458, 0.2065155, -0.1630934, 0.0804516, -0.1999211, 0.0715423, 0.1020874, -0.0994706, 0.0984269, -0.0178563, 0.0775162, 0.0885335, 0.0340338, 0.1005764, 0.1190967, 0.0715478, 0.1342000, 0.0657133, 0.1191710, 0.1684025, 0.1132728, 0.0920322, -0.0332687, 0.1881246, -0.0136231, 0.0610609, 0.1365692, 0.1369737, -0.0021956, 0.0452895, 0.2337901, 0.1041967, 0.1365063, 0.1518371, 0.1537924, 0.0402328, 0.0397852, 0.0697837, 0.1470444, 0.1215085, -0.0165455, 0.0443658, -0.0341164, -0.0451748, -0.1102671, 0.0157457, -0.0362916, 0.1128963, 0.0739777, -0.0428043, 0.1946885, 0.1759533, 0.0171101, 0.1586176, -0.1156489, 0.0754449, 0.0120466, 0.0542424, 0.0646745, 0.0480186, 0.0306618, 0.0331352, -0.1136989, 0.0599178, 0.0933870, 0.0366716, 0.0304879, 0.0584129, -0.0275580, -0.0237591, 0.0004826, 0.1117926, -0.0753477, 0.0113351, -0.0016279, -0.0698601, -0.1979742, -0.0215573, -0.0187232, 0.0802392, -0.0776412, 0.0478428, 0.0451057, -0.1030381, -0.0075960, 0.0787644, -0.0335905, 0.0792335, 0.0386466, -0.1335550, -0.0273603, 0.1545477, 0.2032466, 0.1525761, -0.0057780, 0.0911725, 0.1106340, 0.1333348, 0.0263155, 0.1491454, -0.0030731, 0.0508998, -0.0454749, -0.0670761, -0.0395690, -0.1287903, 0.0599894, 0.1387022, 0.0682064, 0.0770428, 0.0410919, 0.1196038, -0.0293237, 0.0930077, -0.1292014, 0.1584452, -0.0003068, 0.1098755, 0.1524462, -0.0833643, 0.1180828, 0.0810154, -0.0582036, 0.2908887, 0.0917694, -0.2195216, 0.3066523, -0.1254606, 0.2070353, -0.0050783, 0.0850402, -0.0006631, -0.0337750, -0.0604537, 0.1727322, 0.1866926, 0.3555872, 0.1740334, -0.0163356, 0.0401354, 0.2542800, 0.0976098, 0.0011623, 0.4140003, 0.0839449, 0.0974845, 0.2088702, 0.0944115, -0.0987225, 0.0537797, 0.0580811, 0.3601962, 0.1437410, -0.1338037, 0.0905681, 0.1315982, 0.1472212, -0.0144877, -0.0814132, -0.1446063, 0.0164877, 0.0446049, -0.0457486, 0.0151816, -0.0240154, 0.0281498, 0.0727869, 0.0295925, 0.1441139, 0.0566054, 0.1812939, 0.0288403, -0.0007674, 0.0205842, -0.0744104, 0.0671583, -0.0123902, 0.0560656, 0.0396196, 0.0349231, 0.0584414, 0.1169368, -0.0691017, 0.1053287, -0.0138537, 0.0318426, 0.0777090, -0.0094592, -0.0280363, 0.0330309, 0.0484112, 0.0286095, -0.0196183, -0.0631392, 0.0115769, -0.0299093, -0.0286379, -0.0642017, -0.0478327, 0.0971593, 0.2988388, 0.1123401, 0.1377082, -0.1699653, -0.0132192, 0.2047980, -0.2312870, 0.1449994, 0.2710546, -0.1206847, 0.3290255, 0.0832823, -0.2269367, 0.1646780, -0.3424213, 0.2971482, -0.2135608, 0.0045818, -0.0810480, 0.1589883, 0.0971462, 0.2371707, -0.3482259, -0.1915335, -0.2372537, 0.0784005, -0.0076515, -0.2093208, 0.3220437, -0.1148663, 0.4068564, 0.5280769, -0.2922359, 0.4995721, 0.4685331, -0.2902454, -0.0991061, 0.0470047, 0.0082595, -0.3626631, 0.1861437, 0.0205417, 0.0411182, -0.0119296, 0.1631855, 0.0610599, 0.0963765, -0.0399908, 0.2670339, 0.1461879, 0.5319846, 0.0861575, -0.2867419, -0.1794652, -0.1286831, 0.2969329, -0.1845021, -0.0360627, -0.0868371, 0.0578455, 0.2365831, 0.5204930, -0.0969970, 0.1421475, 0.0028103, 0.0345658, 0.1853835, -0.2463242, 0.2720861, 0.0406451, 0.2420362, 0.2820660, -0.4872227, 0.2402731, 0.1409660, -0.3055190, 0.1126225, -0.1107423, 0.2028195, 0.0044556, 0.1192515, -0.1872885, -0.0593440, 0.0694387, 0.2778220, 0.0738573, 0.1730137, -0.0235084, -0.0226290, 0.1208583, 0.2414604, 0.2625857, -0.0777585, 0.0625416, -0.2775479, 0.2042824, 0.1402638, -0.3353551, 0.1058312, 0.2849213, -0.1123308, 0.3297330, -0.3040713, 0.1138975, 0.1640606, -0.2766732, -0.1218511, -0.2780320, 0.2298046, 0.3089083, 0.2807366, 0.2669269, -0.1564563, 0.0361017, 0.1640959, -0.3081996, 0.3864939, 0.1204457, -0.0064470, -0.1720168, 0.1377919, 0.0389443, 0.0387559, 0.3915120, -0.0673484, -0.3652236, 0.4399929, -0.2822309, 0.1227458, -0.0846429, 0.0017237, -0.2612666, -0.2117972, -0.3218226, 0.2561002, 0.0395349, 0.3581111, 0.1127926, -0.0902267, 0.0139275, 0.5953592, 0.0173768, 0.1571457, 0.4539924, -0.0428054, 0.1543698, 0.3787564, 0.1119394, -0.3077905, 0.0058093, 0.0002015, 0.5401369, 0.1264900, -0.2504345, 0.1431586, 0.2001760, 0.0939960, -0.0928359, -0.0007854, -0.0206173, -0.1793898, -0.0331424, -0.0261673, -0.0626082, -0.0347157, -0.1982937, -0.0025181, -0.1343691, -0.0438384, 0.1203210, -0.0334684, -0.0114504, -0.0070930, -0.0305072, -0.1439430, -0.0092754, 0.0816464, -0.0296698, -0.0908308, -0.0610403, -0.0426432, -0.0298215, -0.0571973, -0.0593298, 0.0780718, -0.1269794, -0.0120518, 0.0536390, -0.1720854, -0.0554136, -0.0958712, -0.0659067, -0.0591785, -0.3273630, -0.2150855, 0.0320434, 0.0425613, 0.0680399, -0.0068045, 0.0816254, 0.0098201, 0.0773557, 0.0092134, 0.0788436, -0.0206523, 0.2284243, 0.1248810, 0.0468098, -0.0033982, 0.0746472, 0.1379817, 0.1328840, 0.1498692, 0.0926257, 0.0198589, -0.0186346, 0.0730619, 0.0817366, 0.1527085, 0.1336768, -0.0111482, 0.1012520, 0.0077574, 0.2058170, 0.1137218, -0.0904029, 0.0804215, 0.0676954, 0.0375735, 0.1007465, 0.1347875, -0.0044481, 0.1047996, 0.0464477, 0.1082312, -0.0370181, 0.1156095, -0.0101961, -0.0951231, -0.1245917, -0.0146419, 0.0350655, 0.0190507, 0.1160146, -0.1145869, 0.0584809, 0.1026273, 0.0302292, 0.1817964, 0.0312560, 0.1017510, -0.0723604, -0.0162015, -0.0449103, -0.0903824, 0.0710624, 0.0239840, 0.1112238, 0.0095890, -0.0250868, 0.1784145, 0.1333169, -0.0031945, 0.2363924, -0.0768384, 0.1049030, 0.1184461, -0.0202729, 0.0500306, 0.0227964, 0.0287824, 0.0365443, -0.0526370, -0.0277013, -0.0221650, -0.0647777, 0.0276641, -0.1234723, 0.0003602, 0.1125184, -0.0309323, 0.0038955, 0.0854129, -0.1446476, -0.1418601, 0.0466625, -0.0406221, 0.1407910, -0.0435257, -0.2484493, -0.0818548, 0.1223912, 0.1198404, 0.1447160, -0.2121882, -0.0109377, 0.1367334, 0.0983764, 0.1492435, 0.1676107, -0.1429542, -0.0385397, -0.1670504, -0.0533673, 0.0222603, -0.1336903, 0.0329160, 0.1250223, -0.0213260, 0.1042041, 0.1240109, -0.1439433, 0.0345146, -0.0279982, -0.1231711, 0.0193808, 0.0208832, 0.0447722, 0.0919719, -0.4348463, 0.1099889, 0.0632045, -0.3597309, 0.4088650, 0.0772387, -0.3482806, 0.4989928, -0.3869887, 0.2033656, 0.1167869, 0.1103677, -0.1527099, -0.2033854, -0.3511736, 0.2562292, 0.1209433, 0.3148631, -0.0190871, -0.0683114, 0.0245654, 0.5398988, 0.2213929, 0.0931492, 0.5172530, 0.1312681, 0.0261958, 0.3688700, 0.0605160, -0.2904999, -0.0079193, 0.0843430, 0.4442514, 0.0763460, -0.3647243, 0.2077738, 0.1233260, 0.1267418, -0.0262182, 0.0056518, -0.0540471, -0.0747336, 0.0305997, 0.0132580, -0.0263063, -0.0130357, -0.0224539, 0.0848881, 0.1116477, -0.0069392, 0.0296429, 0.0644631, 0.0289449, 0.1008526, 0.0470207, -0.1180701, -0.0628582, 0.1165816, 0.0700980, 0.0530869, 0.0014300, -0.0167940, 0.0637096, -0.0424711, 0.0506619, 0.0543348, -0.0044639, 0.0692845, 0.0555420, -0.0466852, 0.0735248, -0.0010837, -0.0067833, -0.0126671, -0.2744603, -0.0959141, 0.0065633, 0.0483506, 0.1670499, -0.1798349, -0.0895519, 0.4610194, 0.1473142, 0.1101686, -0.1160855, -0.1250468, 0.1256181, -0.1395406, 0.2140544, 0.3283436, -0.0343973, 0.4608465, 0.0048235, -0.2868685, -0.1009265, -0.0902560, 0.3340625, -0.2591005, 0.1809836, -0.1717378, -0.0007409, 0.3477389, 0.2936395, 0.0520996, -0.0126017, -0.2846230, 0.2605443, 0.2433962, -0.3256636, 0.2151349, -0.2564901, 0.4963197, 0.5440398, -0.4152400, 0.4997355, 0.4752181, -0.3805833, -0.2624646, 0.0062936, -0.0722787, -0.1942495, 0.3576794, 0.0630903, 0.0994782, 0.1098451, 0.0072910, 0.0796826, -0.0021496, 0.0999271, 0.1884199, 0.0852991, 0.4703493, -0.0832146, -0.3796009, -0.1950777, -0.0091594, 0.2048724, -0.1867015, 0.1108488, 0.0440779, -0.1571422, 0.3207128, 0.3995754, 0.1055528, 0.1145609, -0.1554625, 0.1925780, 0.3595253, -0.2505255, 0.2506922, -0.1956612, 0.3429440, 0.3707172, -0.2826610, 0.3094282, 0.4142587, -0.4275095, -0.0746859, 0.0171100, 0.0730404, 0.0907141, 0.0530252, 0.1571360, -0.2866067, 0.0701592, 0.0741167, 0.1158678, 0.1641131, -0.1979062, 0.0089943, 0.2291482, 0.2080244, 0.2089589, -0.1591100, 0.0922381, -0.1858249, 0.0638479, 0.1372337, -0.2184754, 0.0673437, 0.2462169, -0.0291914, 0.1187766, -0.3088259, 0.1582020, 0.0978181, -0.2196802, -0.1024041, -0.2211508, 0.0328913, -0.0025391, 0.1623135, 0.3371685, -0.1668054, 0.1798512, 0.0857301, -0.3221559, 0.1036849, 0.0450271, 0.0330641, -0.1593151, 0.0970069, 0.0314226, -0.0838247, 0.3480336, 0.0093310, -0.2095730, 0.4082309, -0.2890306, 0.1482041, 0.0406616, 0.0654208, -0.2467554, -0.2629621, -0.2075677, 0.1726722, 0.0361294, 0.2424699, 0.0107898, -0.0774453, 0.0280541, 0.4881683, 0.0795325, 0.1601608, 0.3226340, 0.0239233, 0.1017481, 0.1230806, 0.0155105, -0.1420681, -0.0847912, -0.0521275, 0.5138692, 0.0287008, -0.1563174, 0.1453847, 0.1581772, 0.1109874, -0.0786642, -0.0386410, 0.0033360, -0.1875314, -0.0201762, -0.0139397, -0.0480480, -0.0153843, -0.0082193, -0.0093948, -0.0503378, -0.0079735, -0.0902627, -0.0052990, -0.0042091, -0.0118325, 0.0242042, -0.1516264, 0.0152666, 0.0049824, -0.0222649, -0.0003852, -0.0517072, -0.1053946, -0.0462713, -0.0552258, -0.0131878, 0.0373184, -0.1445853, -0.0903352, -0.0176579, -0.0330238, -0.0212356, -0.0624281, -0.0664068, -0.0359990, -0.1200625, -0.2234045, -0.0293671, 0.0096817, -0.0494740, 0.0455239, 0.1050853, 0.0932988, 0.0278060, 0.0696514, 0.0581872, 0.1377768, 0.2254261, 0.0643620, 0.0604248, 0.1024217, -0.0283198, 0.1473244, 0.1191478, 0.0137482, 0.0931584, -0.0263561, 0.1296489, 0.1473851, 0.0396393, 0.1347998, 0.1341286, -0.0556399, 0.2353858, -0.0945846, 0.1330387, 0.0062254, -0.0711529, -0.0131235, -0.0231224, 0.1850649, 0.0694537, 0.1089947, 0.1317658, -0.0423838, 0.1888186, 0.0578817, -0.1096831, 0.1125194, -0.0697554, 0.0320127, -0.0033540, -0.0228994, -0.0394308, -0.0098335, 0.1560363, 0.0412658, -0.0220824, 0.1112884, -0.0330003, 0.0060461, 0.0856883, 0.0153469, -0.0646200, 0.0114129, 0.0033960, -0.0359980, 0.0569534, 0.1244714, -0.0266926, 0.0547998, -0.0001601, 0.0495224, 0.0655212, 0.0014434, 0.1786877, 0.1298510, -0.0723743, -0.0326288, 0.0136847, 0.0345846, 0.0079532, -0.0733898, 0.0528793, 0.0567884, -0.1049796, -0.0524682, -0.0304216, 0.0844451, -0.0069447, -0.0441413, 0.1195807, 0.1014019, 0.0531755, 0.1103237, -0.1843649, -0.0959473, 0.1252143, -0.0735665, 0.1474120, -0.0677915, -0.2295136, -0.0749176, 0.0662781, 0.1147408, 0.1604169, -0.1198273, 0.0749383, 0.0720142, 0.0603380, 0.1216034, 0.1956450, -0.1545039, -0.0273734, -0.1295917, -0.0652463, -0.1011261, -0.0770636, 0.0560220, 0.0788038, 0.0569335, 0.0809412, 0.1531903, -0.0407972, 0.0678087, 0.0702092, 0.0907715, -0.0203202, 0.0289396, 0.0330042, -0.0050513, -0.4135262, 0.1503883, 0.0314686, -0.3259718, 0.5480291, 0.0958754, -0.3103179, 0.6311474, -0.5105738, 0.1450622, 0.1511797, 0.0748356, -0.1738697, -0.2549805, -0.3210726, 0.2997277, 0.0652582, 0.4610186, 0.0255987, -0.0242815, 0.1208379, 0.5384480, 0.1249555, 0.1187448, 0.6162794, 0.1376296, 0.0570522, 0.4477145, 0.0880153, -0.3639096, 0.0384975, 0.0339766, 0.5557261, 0.1482300, -0.3677889, 0.1398166, 0.1675832, 0.2520676, -0.0620774, 0.0003876, 0.0798439, -0.0186235, 0.0195365, 0.0829075, -0.0563909, -0.0604337, 0.0578927, 0.0111378, 0.0726417, -0.0687089, -0.1466314, 0.0096214, 0.0627054, 0.0558374, 0.1097583, -0.0826037, -0.0097801, 0.1264265, 0.0664511, 0.1029697, 0.0667174, -0.0946209, 0.0511102, -0.0397789, -0.0243915, 0.0120654, -0.0442428, 0.0355216, 0.0550433, 0.0396268, 0.0684592, 0.0761173, -0.0899202, -0.0163637, -0.0902096, -0.0300818, -0.0419956, 0.0616485, 0.2000114, 0.1470053, -0.0942704, 0.4905666, 0.0034496, 0.0499601, 0.0853319, 0.1431602, 0.1093294, -0.1093214, 0.2704048, 0.0399934, 0.1675333, 0.1078180, 0.1364946, -0.0329902, -0.1668003, 0.2285554, 0.1298034, -0.5797328, 0.0915425, -0.0580101, -0.0086998, 0.4742438, 0.3611352, 0.2338131, 0.0030657, -0.0300428, 0.3120054, 0.3361648, -0.4228017, 0.1458790, -0.1154589, 0.4439107, 0.2721490, -0.4811943, 0.2148338, 0.5154147, -0.3428074, -0.3314411, 0.0004704, 0.1097581, -0.0852659, 0.2593429, -0.1459782, 0.1024382, 0.1251035, 0.1880468, -0.0350232, 0.0568270, 0.1716027, -0.1070591, 0.1912267, -0.1972643, 0.1795149, 0.1198986, -0.1177282, 0.2570571, -0.0103784, -0.0244696, -0.0541506, -0.0299530, 0.1688226, 0.2448757, 0.2278139, 0.1082779, -0.0828682, -0.0002057, 0.0870182, 0.2437141, -0.1044253, -0.0420522, 0.1890922, 0.2290731, 0.0753013, -0.0172008, 0.0177787, 0.2687474, 0.0226694, 0.1100518, 0.2586488, -0.0064749, 0.2403210, 0.3227348, 0.1764175, -0.1541852, -0.0063471, -0.0429116, 0.2597132, 0.0126134, -0.1716055, 0.0683106, 0.1212996, -0.0033971, 0.3108877, -0.2539722, 0.1911371, -0.0106891, 0.0832401, 0.0694694, -0.2050167, -0.1166155, 0.2731226, -0.0453170, -0.0639554, -0.1648361, -0.0376571, -0.0174075, -0.2267740, -0.2536811, -0.1399457, 0.0081388, -0.0978235, 0.2988227, 0.3290609, -0.0821695, 0.2197722, 0.2689217, -0.2177416, 0.0184580, 0.0866096, 0.0520744, 0.1269411, 0.0905461, 0.0525305, -0.1162458, 0.1787702, 0.0213470, 0.1097693, 0.0771304, 0.1917312, 0.0642247, 0.0083258, 0.0575582, -0.0323757, -0.0002498, 0.1241412, 0.0944091, -0.0659979, 0.0251306, -0.0150423, 0.1378819, 0.0139196, 0.0455451, 0.0638838, 0.0967420, 0.2895013, 0.0764569, 0.0490152, -0.0037655, -0.0737846, 0.1537126, -0.0085731, -0.0168600, 0.0950593, 0.0341970, 0.0538008, 0.0857948, -0.0844133, 0.0901934, -0.0615327, -0.0501299, 0.0004603, -0.1675837, -0.0238916, 0.0064905, -0.0196238, -0.0175939, 0.0042022, 0.0265018, -0.0033317, -0.0033919, -0.0244207, -0.0158069, -0.0140298, 0.0066645, 0.0289326, -0.0948613, -0.0378558, 0.0650318, -0.0090887, -0.0144563, -0.0144331, -0.1070487, -0.0833646, -0.0234573, 0.0042749, -0.0096552, -0.0904427, -0.0761769, 0.0104986, -0.0315157, 0.0119706, -0.0763328, -0.0547257, 0.0153663, -0.0890125, -0.1935240, 0.0115405, 0.0110074, 0.1994217, 0.0472024, 0.0695903, 0.0774291, 0.1151131, 0.0432803, -0.0242709, 0.1525495, 0.2583062, 0.0192257, 0.1411268, -0.0580435, 0.1413283, 0.0678855, 0.1869601, 0.0133453, 0.0823341, 0.0571003, -0.0429139, -0.0383771, -0.0352478, 0.0556470, 0.1028171, -0.0368332, 0.0830408, -0.0009274, 0.0538294, 0.0207160, 0.0881187, 0.0221356, -0.1131435, 0.1756865, 0.0644833, 0.1141767, 0.1311429, -0.1245274, 0.1681888, 0.1515808, -0.0965803, 0.0330318, -0.0537257, 0.0063922, -0.0203359, 0.0084222, 0.0210339, -0.0074029, 0.0867490, 0.0898741, 0.0200370, 0.0796753, -0.0527399, -0.0308679, 0.0539219, 0.0144492, -0.0123425, -0.0506877, 0.0064752, 0.0434674, -0.0068482, 0.0062393, -0.0569170, 0.0490925, 0.0418604, 0.0549713, 0.0839146, 0.0007872, 0.0717217, -0.0055607, -0.0618955, -0.0093869, -0.0866237, 0.0037499, 0.0114391, -0.0236769, 0.0694976, -0.0025127, 0.0193551, 0.0034353, -0.0410780, 0.0623858, 0.1467549, -0.0581024, 0.0022270, 0.1643768, 0.0940395, 0.0492144, -0.2167602, -0.0781478, 0.0481818, -0.2041931, 0.1334460, -0.0910817, -0.0282759, -0.0467013, 0.1382554, -0.0139197, -0.0201999, -0.0289488, 0.0136933, -0.3611299, 0.0422723, -0.0979542, 0.0893514, -0.0189472, 0.0034756, -0.1276010, -0.2265957, -0.1967098, 0.0530469, 0.0549864, -0.0425771, -0.0176808, -0.0819626, 0.1810920, 0.0314586, -0.2606430, 0.1520295, 0.1224468, -0.1269563, -0.3914556, 0.0126192, 0.0388878, -0.1536678, 0.1307151, -0.0333963, -0.1963573, 0.2391461, 0.0510882, -0.1244044, 0.6535830, -0.3132107, -0.0356444, 0.0621204, 0.0189536, -0.0936341, -0.1144304, -0.1482112, 0.2745925, -0.1950228, 0.3562416, -0.0470132, 0.1122989, 0.1577906, 0.2822900, 0.0901616, 0.0670202, 0.4836394, 0.0463826, -0.0267953, 0.3264292, 0.0769695, -0.1496516, 0.1883902, 0.0669077, 0.2420239, 0.2662615, -0.2848703, 0.1632433, 0.1084637, 0.1958614, -0.1713856, -0.0367995, 0.0804756, -0.0904012, -0.1397588, 0.0827918, -0.0047375, 0.0014405, 0.0177971, 0.0363677, -0.0137240, -0.1662420, -0.2101651, -0.2427445, 0.0142377, 0.0423325, 0.0754040, -0.0134342, -0.0590121, 0.1960151, -0.0424521, 0.1604633, 0.1816481, -0.2106862, -0.0533549, -0.0679546, -0.0263445, 0.0347857, -0.1583365, -0.0811618, 0.0298240, -0.0067292, 0.1648360, -0.0307215, -0.2227040, 0.1197521, -0.1035899, -0.1814564, 0.0397525, 0.1881869, 0.1316010, 0.1821142, -0.3089069, 0.3959805, -0.1435375, 0.1739319, 0.0588043, 0.0842825, -0.1088218, -0.0825999, 0.3018261, 0.1202060, 0.1430113, 0.2633570, 0.0728890, 0.0347470, -0.3516921, 0.0818656, 0.1959192, -0.5080383, 0.1885163, -0.0920216, -0.2201515, 0.4812946, 0.6748853, 0.0529066, -0.1106730, -0.0490377, 0.3011606, 0.5634972, -0.3706664, 0.1174299, -0.1708799, 0.4095572, 0.1231601, -0.5208338, 0.1996432, 0.4552335, -0.3266910, -0.4174153, -0.1806655, -0.1082678, -0.1451999, 0.3187599, -0.2830610, 0.2352955, -0.0283603, 0.1084741, -0.0265265, 0.1079030, 0.0672217, -0.1118049, -0.0436337, -0.1089004, 0.0233533, -0.0555052, -0.1522012, 0.2657837, -0.0022320, -0.1201643, -0.0660707, 0.0608125, 0.1769071, 0.3046165, 0.2860748, 0.0093204, -0.1394739, -0.2369946, 0.1139905, 0.2547652, -0.1476028, 0.1913657, 0.2166635, 0.2136690, 0.1017285, -0.0474752, 0.1861652, 0.3043762, 0.0669261, 0.1609646, 0.1924178, 0.3476614, 0.2059374, 0.1994013, 0.1066410, -0.2226407, 0.0764344, 0.1357722, 0.1271626, -0.1132323, -0.0207320, 0.0857615, 0.2327636, -0.0511855, 0.2941071, 0.0694664, 0.1466394, 0.0365074, 0.0123158, -0.0270268, -0.2668838, -0.1117884, 0.1189766, -0.0451015, -0.0131749, -0.0649833, -0.0318389, 0.3210017, -0.1159365, -0.2893160, -0.0842190, 0.0168760, -0.1811531, 0.1173313, 0.0573206, -0.0907512, 0.0467859, 0.1307873, -0.1736083, 0.0300362, 0.2441764, 0.0959904, 0.3602654, -0.0392414, 0.2707216, -0.1323256, 0.1836012, -0.0685958, 0.2520206, -0.3150762, 0.4600709, 0.2477052, 0.0277592, 0.2292247, -0.0626135, 0.0382561, 0.4754758, 0.2013005, -0.1210555, -0.1796898, 0.0886838, 0.4515303, -0.0031118, -0.3954125, 0.0201857, 0.2278536, 0.1150784, 0.0132730, 0.3961376, -0.2114812, -0.2923396, 0.3170035, 0.0209467, -0.0087296, -0.3419432, 0.1010870, 0.2535166, 0.0495971, -0.3713143, -0.2035313, -0.0384197, -0.0200751, -0.0147901, -0.1242846, -0.0278375, 0.0158010, -0.0736867, -0.0093337, -0.0126296, 0.0509095, 0.0002592, -0.0168833, -0.0207235, -0.0091469, -0.0018393, 0.0100385, 0.0053239, -0.0930819, -0.0164734, 0.0433115, 0.0057904, 0.0144194, -0.0065903, -0.0465914, -0.0417752, -0.0507010, 0.0033431, -0.0178903, -0.0741656, -0.0096143, 0.0090940, -0.0068679, 0.0397115, -0.0400352, -0.0092315, 0.0021931, -0.0499780, -0.1192883, 0.0184476, 0.0565002, 0.1751693, 0.0929120, -0.1199987, 0.4384114, -0.0963694, 0.2170753, -0.1101168, 0.0904524, -0.0552322, -0.3198740, 0.4677754, 0.0553308, 0.0313105, 0.0370699, 0.1466268, 0.0718206, -0.2228911, 0.1285834, 0.0917645, -0.4633000, 0.1460574, -0.2479379, -0.1882592, 0.3790498, 0.3800100, 0.0628748, -0.3131038, -0.0414280, 0.5170066, 0.4022788, -0.1901032, 0.1411358, -0.1158994, 0.3465876, 0.0705636, -0.3367940, 0.3027516, 0.5119032, -0.2451963, -0.4542469, 0.0808453, -0.0614597, -0.0413901, -0.0335970, 0.0390416, -0.0379898, -0.0083859, 0.0439592, -0.0258952, 0.0445551, -0.0682419, -0.0735027, 0.0076763, 0.0364795, 0.0248987, -0.0103617, -0.0210973, 0.0169331, -0.0955083, 0.0071601, -0.0168643, -0.0413959, -0.0260602, 0.0339191, -0.0133389, 0.0236142, -0.0304398, -0.0294362, 0.0296792, -0.0293348, 0.0078051, -0.1003741, -0.0180513, -0.0013882, 0.0342466, -0.0382750, -0.0095789, -0.0093808, 0.0297263, -0.0258160, 0.1066149, 0.0157146, -0.0778597, 0.1146689, 0.1002938, 0.0747283, -0.1028173, -0.1160688, -0.0767470, -0.1252600, 0.1296500, 0.1071227, -0.0268256, 0.1879564, 0.0261011, -0.0248217, -0.1156650, -0.0338838, 0.1403657, -0.3047616, 0.0862696, -0.2496414, -0.0815321, 0.1764704, 0.1561274, 0.0868743, -0.0863293, -0.1934650, 0.1247127, 0.1497594, -0.0230985, -0.1109613, -0.3086534, 0.2145442, 0.2073096, -0.2074544, 0.0536289, 0.1492158, -0.0408073, -0.5138635, 0.0571957, 0.1485211, 0.2665842, 0.0501734, 0.0605996, -0.1626574, 0.1604993, 0.2141857, 0.2592976, -0.0027869, 0.1038099, -0.0061284, 0.1237531, -0.0443079, 0.0501788, 0.0265911, 0.2534986, 0.2712050, -0.2350744, 0.0291800, -0.1514284, 0.3083934, 0.1160863, -0.1378195, 0.1184853, 0.0276900, 0.0871537, 0.2583148, 0.0981192, -0.2044443, -0.0579285, 0.2971105, 0.1796418, -0.0073709, -0.0692912, 0.1374399, 0.1165554, 0.2305020, -0.1587619, 0.2723843, -0.2098752, 0.0573040, 0.0493372, -0.0885682, -0.1332305, 0.1423364, -0.1498225, 0.0747521, 0.0759700, 0.1217693, 0.0632226, -0.0667142, -0.2266445, -0.1829161, 0.0926449, 0.1018207, 0.0879550, 0.0585019, 0.0013461, 0.2011085, -0.0386637, 0.1102160, 0.1869079, -0.1922160, -0.1257148, -0.1763502, -0.1708822, 0.1077505, -0.1809691, -0.0300265, 0.0505575, 0.1738379, 0.2371485, -0.0685698, -0.1207188, 0.0888228, -0.0251617, -0.1699377, 0.0028815, 0.2721141, -0.1063469, -0.0736812, -0.4974651, 0.2279645, -0.1206848, 0.4253391, -0.1026484, 0.0741363, -0.0452709, -0.1385125, 0.3695145, 0.2328191, 0.0735466, 0.6263177, -0.1106671, -0.1651407, -0.4640736, -0.2949940, 0.3592645, -0.2621064, 0.3326749, -0.0544041, -0.2471756, 0.2760742, 0.6528785, -0.1672275, -0.0261236, -0.1581771, 0.3662385, 0.5918167, -0.2409606, 0.2983925, -0.1848152, 0.4294698, 0.2855980, -0.5080020, 0.2778952, 0.3621129, -0.3521821, -0.2790044, -0.2197759, -0.2181816, -0.2349196, 0.1087736, -0.1407121, 0.4367005, -0.0689837, 0.2414292, 0.0942215, 0.2318544, 0.0617228, -0.0664750, -0.1355433, -0.0460376, 0.1885927, -0.0645974, -0.1862452, 0.3130642, 0.0336972, -0.1248837, 0.0248847, 0.0827793, 0.3094518, -0.0179783, 0.1001004, -0.0171388, -0.0821780, -0.1905898, 0.0072193, 0.0938679, -0.1323628, 0.3363983, 0.3399644, 0.0805869, -0.0503485, 0.0676781, 0.2752511, 0.0536305, 0.2456452, 0.2513930, 0.0919384, 0.0975638, -0.0046983, 0.0640953, 0.0622496, -0.2134320, 0.0418636, 0.0626000, 0.2378218, -0.1208277, 0.0786469, 0.2416392, 0.1477518, 0.4741964, 0.0796648, -0.0489164, 0.0389413, -0.1137629, 0.0845480, -0.2496997, -0.1137837, -0.0010000, -0.0454555, -0.0710000, 0.2880653, -0.0665800, 0.0937228, 0.0931220, -0.0395217, -0.1108826, -0.2464685, 0.1474290, -0.2462319, 0.1292272, -0.0312384, -0.2201162, 0.1973005, 0.1355663, -0.3934059, -0.0719798, 0.1244239, 0.2023631, 0.3175815, -0.0116908, 0.2055204, -0.0347215, 0.1362875, -0.1627939, 0.3064746, -0.3775910, 0.4612233, 0.2797759, -0.0158131, 0.1501463, -0.0382920, 0.0351412, 0.4572094, 0.1788190, 0.0917754, -0.2197319, 0.1778046, 0.2765217, -0.1117904, -0.4208594, -0.0156075, 0.1899773, 0.0786231, 0.2806242, 0.3124118, -0.3294607, -0.1940268, 0.2839465, -0.1451755, -0.0290803, -0.2683584, 0.0894194, 0.1399142, -0.0093123, -0.2190116, -0.1412721, -0.0330010, -0.0462154, -0.0232713, -0.0569949, -0.0057863, -0.0260294, -0.1016895, -0.0412207, 0.0241314, 0.0218294, 0.0126320, -0.0711363, -0.0755152, 0.0054942, -0.0013701, -0.0112929, 0.0299660, -0.0486918, -0.0173889, 0.0101419, -0.0103205, -0.0146525, -0.0241298, -0.0898063, -0.0199624, -0.0404646, -0.0414285, -0.0224483, -0.0706250, 0.0300935, -0.0106493, -0.0298949, 0.0268925, -0.0222100, -0.0990705, -0.0217283, -0.0285468, -0.1257730, -0.0066312, 0.0155052, 0.1522049, 0.0385619, 0.2307205, 0.1028314, 0.1268349, 0.2701571, -0.0933318, -0.1589596, 0.0951257, 0.0324136, 0.0624760, 0.3874061, -0.3262305, 0.1425928, -0.0532328, -0.0804307, 0.1815013, -0.0919679, 0.2995048, 0.1562904, 0.1312381, 0.1061390, 0.1906346, 0.2112647, -0.0840586, -0.2850819, -0.0844631, -0.0886488, 0.1804273, 0.0529491, -0.0343725, 0.2582644, 0.1425748, 0.1414265, 0.4098138, 0.0856328, 0.4094260, 0.2160042, 0.0725264, 0.0579728, 0.0871873, 0.0001443, 0.0183335, 0.0332817, 0.0672033, -0.0031390, -0.0074000, -0.0546331, -0.0059579, 0.0083861, 0.0147908, -0.0168437, -0.0053377, 0.0407504, 0.0086580, 0.0097273, 0.0283632, -0.0469317, 0.0415080, 0.0501401, 0.0245130, -0.0200011, -0.0295705, 0.0049478, 0.0166394, -0.0207092, 0.0376033, -0.0168778, 0.0627262, 0.0260310, 0.0441398, -0.0834839, -0.0291148, 0.0261337, 0.0609764, -0.0271529, 0.0041843, 0.0180362, 0.0237042, -0.0533476, 0.1003652, 0.1309786, -0.0483867, 0.0364096, 0.1561759, -0.0829215, 0.1002434, 0.0116627, 0.0173754, 0.0622522, 0.0511322, 0.1482428, 0.1950043, 0.3401445, 0.0005724, -0.0292347, -0.0437388, 0.0108489, 0.1975377, -0.0954196, 0.0860496, -0.0626562, -0.1942602, 0.1829966, 0.1815397, 0.0725178, 0.1428082, 0.1067795, 0.0486586, 0.1191973, -0.0147145, -0.0942066, -0.2724214, 0.0515946, 0.1912611, -0.1239907, 0.0793045, 0.0391644, -0.0760982, -0.2634875, 0.3682576, 0.0859377, 0.2345161, 0.2112186, 0.2998402, -0.1388068, 0.1281006, 0.1218131, 0.5181636, -0.2024727, 0.0156062, 0.0818980, 0.1134205, 0.1041523, 0.1693329, -0.0086176, 0.3934056, 0.0868326, -0.0861020, -0.1469483, -0.1295395, 0.1384254, 0.1579932, -0.2651982, -0.0778029, 0.1239410, 0.0132990, 0.0777871, 0.0467952, -0.3538707, -0.1623498, 0.2041722, -0.0213068, 0.1247711, 0.1483202, -0.0464749, 0.4645438, 0.3038452, -0.3164675, 0.0444863, -0.0575711, -0.0136898, -0.0190240, -0.1021003, -0.0011385, 0.1955071, -0.3970118, 0.1167965, 0.1664696, 0.1121326, 0.0026313, -0.1852220, -0.0285514, -0.2733344, 0.3560500, 0.1895644, 0.0911999, 0.0779006, -0.0461686, -0.0882405, -0.0012991, -0.0808129, 0.3391721, -0.3622526, -0.1073313, -0.0749530, -0.2513201, -0.0286114, -0.2231511, -0.1116854, 0.1331037, -0.0142086, 0.1840472, 0.0455690, -0.2703449, -0.1408923, 0.0816676, -0.1141129, 0.1381859, 0.1069678, 0.1006680, -0.0781521, -0.0949109, 0.0787159, 0.0521968, 0.1256442, -0.1038022, 0.0204933, -0.0282639, 0.1828384, 0.2373559, -0.0258177, -0.1203942, 0.1140800, 0.0696011, 0.0625215, 0.0728868, 0.0306527, -0.0453505, -0.0019202, 0.1357486, 0.2689219, 0.0240443, 0.2270088, 0.1567024, 0.0595743, 0.1400940, -0.0268193, 0.0108888, 0.3795638, 0.0828789, -0.0788583, 0.1804249, 0.4004452, 0.1272852, -0.0975064, 0.0691007, 0.2122436, -0.1054861, -0.1607567, 0.0277759, -0.1280569, 0.0269636, -0.0888978, 0.0932449, 0.2017203, -0.1054327, 0.1543622, 0.3284515, 0.1647579, 0.0747022, -0.0258759, 0.0063146, 0.2006258, 0.0939488, 0.0642420, 0.1048628, 0.1364525, -0.0636652, -0.0928193, 0.0544686, 0.1341979, 0.1183528, -0.0831060, -0.0366382, 0.0767121, -0.0278421, -0.0251067, 0.1020584, -0.0103325, -0.0288234, 0.0963015, 0.1671385, -0.0373385, -0.2165584, -0.0691990, 0.1656215, -0.0887564, -0.0325916, 0.0247777, 0.0846544, -0.1046203, 0.1145490, 0.2131162, 0.1889103, 0.0748692, 0.0017371, -0.0692868, 0.3358645, -0.1293322, 0.4714379, 0.2408403, 0.0755061, 0.7831920, 0.1281818, 0.0771533, 0.1604212, -0.1080826, 0.1184970, -0.0728125, 0.2252396, 0.4374176, 0.0124639, -0.0397824, 0.4530437, 0.0658314, 0.2300296, -0.0702217, 0.1837623, 0.0823272, -0.1325050, 0.1879413, 0.1807942, 0.3953682, 0.0867725, -0.1734515, 0.2963832, 0.2190295, -0.5275363, -0.2011368, 0.1088382, -0.0126250, 0.2242710, 0.1535937, 0.0593458, 0.0485970, 0.0243252, 0.0833854, 0.3206502, -0.3279304, 0.2811354, 0.1753653, -0.1561201, 0.2097505, 0.0739568, 0.0534517, 0.3563182, 0.0557078, 0.0325506, -0.1890330, 0.1334808, 0.2167464, 0.0065916, -0.2893002, 0.1032380, 0.0657904, 0.0104213, -0.0374572, 0.1672561, -0.1586616, -0.0880480, 0.4142688, -0.0382136, 0.1144928, -0.1537159, 0.0979753, 0.3183020, 0.1227303, -0.2797606, -0.1695196, 0.0465881, -0.0443621, -0.0860672, -0.0709383, 0.0589871, -0.0036913, -0.0610286, 0.0502912, 0.0472779, -0.0341388, 0.0465347, -0.0480031, -0.0114475, 0.0526775, 0.0669345, 0.0066723, 0.0272468, -0.0855034, -0.1073134, -0.1062993, 0.0170252, -0.0373747, -0.0459504, -0.2028601, 0.0648094, -0.0359135, 0.0098846, 0.0066875, -0.0542800, -0.0146714, -0.0507693, -0.0472546, -0.0207496, -0.0234011, -0.1907020, -0.0890059, 0.0054531, -0.1653658, -0.0718533, -0.1134041, 0.2516937, 0.1196726, 0.3588760, 0.2140131, 0.3244825, -0.0396469, -0.0389662, 0.0371179, 0.1499780, 0.2236769, -0.1928027, 0.1000544, 0.0906281, 0.0223210, 0.3025897, 0.0241231, 0.2916668, -0.1520069, 0.2293301, 0.2248868, 0.0553297, -0.0841220, 0.1741064, -0.0303105, -0.0268581, -0.1598759, -0.0095557, 0.2452289, -0.2756846, -0.1034037, 0.1594044, 0.0006581, -0.1184837, 0.1701616, 0.2688566, -0.0318796, 0.0973513, 0.1421477, 0.1554397, 0.2059351, 0.0724534, -0.0711373, 0.0172192, 0.0547087, 0.0391995, 0.0285420, 0.0214514, 0.0223538, 0.0652986, -0.0064204, 0.0503847, -0.0013499, -0.0322227, 0.0306770, 0.0373024, -0.0152507, 0.0407067, 0.0537323, -0.0634527, -0.0236006, -0.0144830, 0.0510025, -0.0026817, -0.0791094, 0.0952204, 0.0092500, 0.0192566, -0.0833301, 0.0267728, 0.0365224, -0.0222195, 0.0137222, 0.0144680, 0.0481237, -0.0210899, -0.0199296, 0.0369358, -0.0156874, -0.0305373, -0.0409125, 0.0348651, 0.0489496, -0.0415854, 0.0447810, 0.0166361, 0.0426537, 0.0920335, 0.1103149, 0.0420036, -0.0359087, 0.0658759, 0.0561400, 0.0524910, 0.2461255, 0.0747976, -0.0008786, -0.0571616, -0.0721772, 0.2068473, -0.0439886, 0.0183057, -0.0273910, -0.1956877, 0.0558618, 0.2112536, -0.0292147, 0.0594235, 0.0069810, 0.0711564, 0.0704586, -0.0711378, 0.1093285, -0.0991039, 0.0821107, 0.0769653, -0.1124661, 0.1263391, 0.0796445, -0.0950512, -0.0196921, 0.3221885, -0.0248847, 0.2230624, 0.1373910, 0.2750359, -0.0991246, -0.0645010, 0.0360085, 0.3319415, -0.2748961, 0.1055813, 0.0441116, 0.0253308, 0.1857257, 0.1318336, 0.0105254, 0.3962411, -0.0467170, 0.0295718, -0.1215806, 0.0031421, 0.1169323, 0.1679467, -0.0970057, -0.1023344, 0.0627370, 0.0251556, 0.0464199, 0.1181006, -0.0818960, -0.0611394, 0.1192609, -0.0442265, 0.1943934, 0.2394320, -0.1096103, 0.2456082, 0.3405989, -0.3143480, -0.1795442, -0.0833087, 0.0030893, -0.1174655, -0.1450526, -0.0446197, 0.0022211, -0.1227050, 0.0473780, -0.0646364, 0.0005346, 0.0200203, -0.0285478, 0.0617736, 0.0687028, 0.0570864, -0.0160527, -0.0504995, -0.1361750, 0.0151053, 0.0099778, 0.0382737, -0.0697767, 0.0077905, -0.0608993, -0.0104459, -0.0889746, -0.1164314, -0.0103696, -0.0432220, -0.0214681, 0.0307001, 0.0173161, 0.0050087, -0.0527698, -0.0286224, -0.1215084, -0.0437134, -0.2288861, -0.0331029, 0.0146221, -0.0026864, 0.2241103, 0.1953837, 0.1674552, -0.1658006, 0.2416267, -0.1062032, 0.1285445, 0.1027052, -0.1358036, -0.0462326, -0.0155769, -0.0098869, -0.0498505, 0.0524429, 0.1037508, -0.0113547, 0.0949071, 0.1576162, 0.0476510, -0.0102740, -0.2947520, -0.0598238, -0.0545425, -0.1178133, -0.0080228, -0.2530836, 0.0998762, 0.1417874, -0.0627249, -0.0758275, 0.2062505, -0.0905477, -0.0190830, 0.0370357, 0.0358082, 0.2498071, 0.1575051, 0.2565734, 0.1328678, 0.1879598, 0.0292055, 0.0283642, -0.1379514, 0.3222058, -0.1913233, 0.2443041, -0.0050178, 0.0679849, 0.1016677, 0.1511962, 0.0164213, 0.0053454, 0.3648182, 0.1230515, 0.2046283, 0.0836347, 0.1653456, 0.1425128, 0.2641229, 0.3013302, 0.2750333, 0.1017017, 0.0908281, 0.1144869, 0.1640176, 0.3260494, 0.1452681, 0.1229191, 0.1631760, 0.1830950, 0.0805257, 0.1213675, 0.1448772, 0.0795954, 0.1520004, -0.0893272, 0.0114161, -0.0696175, 0.1495796, 0.1551785, 0.1066879, -0.1609744, 0.1288498, 0.0802042, -0.1841685, 0.5991416, -0.0785116, -0.1675892, 0.5992017, -0.1354745, -0.0426798, -0.0568932, -0.0273967, -0.2379935, -0.0425589, -0.1186791, 0.4636391, -0.0536691, 0.5096235, 0.2402264, 0.1855046, 0.0135867, 0.4575522, 0.0567586, 0.1282387, 0.6322478, -0.0065180, 0.1061429, 0.3383338, 0.0720210, -0.1843681, 0.1229748, 0.1136992, 0.4564906, 0.4151947, -0.0965243, 0.2323687, 0.2482786, 0.1243666, 0.1133336, -0.0230323, -0.3216505, 0.0835781, 0.0798696, -0.3053403, 0.4165521, 0.1053860, -0.2015072, 0.6096989, -0.2519154, 0.0411389, 0.1338859, 0.0273263, -0.0110251, -0.1591887, -0.1672491, 0.2123935, 0.0429528, 0.4604957, -0.0771231, -0.0240739, 0.1049104, 0.4384114, 0.1880401, 0.0614208, 0.5837247, 0.0528890, -0.0266782, 0.1995142, 0.0162510, -0.0778056, 0.0650994, 0.0215151, 0.4394090, 0.0284875, -0.1550942, 0.0798885, 0.0430576, 0.1287125, -0.0792140, -0.0363567, -0.1601450, -0.0478834, -0.0030997, 0.0281500, -0.0203277, 0.0984934, -0.1005459, 0.1984915, -0.1632164, -0.1784325, 0.0746087, -0.0407575, 0.2007479, -0.0858410, -0.2329829, 0.0036999, 0.0710610, 0.1230620, -0.1125834, -0.0161373, 0.1371813, 0.1506927, 0.0361896, -0.0541036, 0.0650370, 0.0046743, -0.2090179, 0.2011981, 0.1047939, -0.0669482, 0.2261301, 0.0495058, 0.0769094, -0.0887442, -0.1629572, -0.0631981, 0.0428292, 0.1855581, -0.0346689, 0.1449112, 0.1624257, -0.0837277, 0.0418568, 0.0274392, -0.1957526, -0.1367159, 0.0902876, -0.0834332, 0.1746452, 0.0164768, -0.1128787, -0.0505432, 0.1231580, 0.1125871, 0.2103740, -0.1869104, 0.0156295, 0.0175806, 0.1350886, 0.2188683, 0.1159448, -0.1943038, 0.0208611, -0.1124082, -0.0535327, -0.0096759, -0.1397816, -0.0212330, 0.0951706, 0.1319864, 0.1114678, 0.1783789, -0.0743758, 0.0139321, 0.1253486, -0.1136980, -0.0198630, 0.0060518, -0.1328539, 0.1931229, 0.0485803, -0.1283132, -0.0649556, 0.0189595, -0.1565095, 0.0334692, -0.0826765, 0.0210446, 0.0165446, -0.0576830, 0.1052079, -0.0355089, 0.0985410, 0.0663263, 0.0580203, -0.3104337, 0.1827456, 0.0618886, 0.0482693, -0.1233096, 0.0390197, -0.0574384, 0.0359619, -0.2677861, -0.0792790, 0.1703481, -0.2033022, -0.0168509, 0.0331390, 0.0387186, -0.0542359, -0.0215555, 0.0166664, -0.0581189, -0.0454043, -0.1566454, -0.0233822, 0.0995279, -0.1608906, 0.1316460, 0.1242543, -0.0569359, -0.0783278, 0.2661624, -0.3683412, 0.1543455, 0.0598768, -0.0456924, 0.0386602, -0.0201069, -0.0319946, -0.1479166, 0.1769896, 0.2352724, 0.0836639, 0.0121144, 0.1445604, 0.0293939, 0.0518997, -0.1530436, 0.1266800, -0.2086044, -0.1035847, -0.0321010, -0.2482962, 0.0888532, -0.1140700, -0.0975460, 0.1271202, 0.1708219, 0.0257097, 0.0284604, -0.1045096, -0.0781363, 0.0276988, -0.0310144, 0.2224044, 0.1199587, 0.0554343, -0.0153441, -0.2010548, 0.0429024, 0.0806578, -0.0629874, 0.0555024, 0.0373088, -0.0530086, 0.2337139, -0.0162769, 0.0144244, 0.0786947, 0.0706406, 0.1224032, -0.0135454, -0.0052537, 0.0257387, -0.0005925, 0.1679812, 0.0314911, 0.0470602, 0.1242037, 0.2594190, 0.1702985, -0.0958203, 0.2050693, 0.0877495, -0.0377123, 0.1276651, 0.0466496, -0.0439129, 0.0880544, 0.0113309, 0.1537482, -0.0728617, -0.2123297, -0.0584227, 0.0315954, -0.0133661, -0.0552762, -0.0541618, 0.0464481, -0.1287360, 0.0545000, 0.0961014, -0.0400670, -0.0966791, -0.0062033, 0.0460477, 0.0862605, -0.0022164, -0.0973242, 0.0856203, 0.0298137, 0.0509251, 0.0495826, -0.1342449, 0.0072677, 0.0741507, 0.1188542, 0.0522000, 0.0419188, -0.0872158, 0.0304471, -0.0847600, 0.0618811, -0.0127089, -0.0703449, -0.0094747, 0.0449082, -0.0840152, 0.1096401, 0.0327092, -0.1068498, -0.0257348, -0.2257089, -0.2500864, -0.0186634, -0.0192221, 0.2105472, -0.0859121, 0.1908251, 0.3843774, 0.1468824, 0.1081790, -0.2811216, -0.0192613, 0.2981529, -0.2238428, -0.0123710, 0.0986557, -0.1380368, 0.1189851, 0.1451598, -0.3355972, 0.0530828, 0.0570462, 0.2230386, -0.2695850, 0.0421720, -0.3239979, 0.1482777, 0.0594661, -0.1235203, -0.0356842, -0.2446515, -0.2577297, 0.1696722, -0.0138806, -0.1499503, 0.1246586, -0.1652778, 0.2904641, 0.4209167, -0.0955572, 0.6100873, 0.3717089, -0.0365663, -0.1395158, 0.0767506, -0.2519256, -0.0368647, 0.3039175, 0.1691742, -0.1381512, 0.1321342, -0.1846714, 0.0476911, 0.0798097, 0.2339923, 0.0369551, -0.1586815, 0.2148515, -0.0070897, -0.0619587, 0.0788525, 0.0011940, 0.0162507, 0.0467682, 0.1697914, 0.3565756, 0.0620357, 0.2040039, 0.2707261, -0.0105153, 0.1961739, -0.2103415, 0.0765967, 0.3171118, 0.0391847, 0.0448951, 0.1045501, 0.3278389, 0.2128997, 0.1943174, 0.0505998, 0.2645461, -0.1785629, -0.0203460, -0.0913919, 0.0857885, 0.0341921, 0.2172760, -0.1071366, -0.1448381, 0.3878433, -0.0642658, -0.1389362, 0.2567745, -0.2984727, -0.0448872, -0.0280497, -0.1387529, -0.2844758, -0.3097162, -0.1500737, 0.2835856, 0.0347555, 0.3119032, -0.1764193, 0.0857014, 0.1062693, 0.3672079, 0.0863678, -0.0879859, 0.2642325, 0.0496926, -0.3249004, 0.0911662, -0.0972484, -0.1964113, -0.0157160, 0.1128995, 0.4125881, 0.1635762, -0.0560345, 0.1992682, -0.0206690, 0.2305799, 0.1221883, -0.0082116, -0.3382972, 0.1024877, -0.0160145, -0.4319973, 0.5524691, 0.1513111, -0.2170501, 0.3818114, -0.5451081, 0.0759609, 0.1765633, 0.0912237, -0.1622235, -0.3491019, -0.3417107, 0.2440195, 0.0278009, 0.2022795, -0.1811278, -0.0616181, -0.0075408, 0.5478415, 0.1753195, 0.2198563, 0.5077182, 0.0743916, -0.0254130, 0.1321325, -0.0648419, -0.1175653, -0.0262132, -0.1199089, 0.3464497, -0.0764980, -0.4351294, 0.1134734, 0.0436404, 0.0908339, -0.1256177, -0.0237269, -0.1159206, -0.0121764, -0.1304316, 0.0594921, -0.0391829, 0.0186382, -0.2029642, 0.0679089, -0.1403684, -0.0994834, -0.1456499, -0.1224966, -0.1432206, -0.0436422, -0.1778080, 0.0192312, 0.0296480, 0.0338924, -0.0430954, -0.1258576, -0.0400376, 0.1483805, -0.0768703, 0.1072767, -0.0594078, -0.0235436, -0.0500668, 0.1896669, 0.0200122, -0.1244803, 0.1029991, -0.0683164, -0.0706017, 0.0493115, -0.1188099, -0.0203394, 0.1192319, 0.0799467, -0.1554596, 0.0310403, 0.0680020, -0.1035245, -0.0240219, 0.1251769, -0.1658268, -0.0475126, 0.1850318, -0.0407326, 0.1776800, 0.0565171, -0.2836691, 0.0331621, 0.0700190, 0.1082582, 0.1473857, -0.1506450, 0.1255077, 0.0920704, 0.0834126, 0.0524614, 0.0928745, -0.2889499, 0.0243712, -0.1208974, -0.0503689, 0.0222295, -0.1130742, -0.0711102, 0.0486675, 0.2141496, 0.0705790, 0.0731339, -0.0991558, -0.0061539, 0.0968491, -0.0891670, 0.0190885, 0.1047643, -0.1846271, 0.0098500, -0.0169917, -0.1714063, 0.0281997, 0.0382620, 0.0252183, -0.0505869, 0.0365964, 0.1334455, -0.0656190, 0.0665896, -0.0430537, 0.2285143, -0.0357428, -0.0586245, 0.1316602, -0.2677960, 0.1617613, 0.1582134, -0.0523062, 0.0597175, 0.1538630, -0.0490622, 0.2107692, -0.2175450, 0.0896969, 0.0711305, -0.2353833, -0.0907738, 0.0387738, 0.0095953, 0.1421679, 0.0330925, 0.1484927, -0.1143543, -0.1395476, -0.2725442, -0.0630374, 0.1131137, -0.2228918, 0.1507777, 0.1192001, 0.0072301, -0.0255048, 0.1816597, -0.1765456, 0.0335548, 0.0676885, -0.0262520, 0.2002735, 0.0416730, -0.2692401, -0.1279450, 0.0770853, 0.1197400, 0.1562399, -0.1180852, 0.2226943, 0.0860561, 0.1698504, -0.0727434, 0.1648474, -0.1336323, -0.0754054, -0.1378912, -0.1579282, 0.0732771, 0.0124626, 0.0060216, 0.1051987, 0.1162878, 0.0149246, 0.0691232, -0.0554199, 0.0171287, 0.0435259, 0.0213232, 0.0847165, 0.0892196, -0.0093982, -0.0147665, -0.2878943, 0.0481997, 0.0048496, -0.2349518, 0.0528008, -0.0722859, -0.0843332, 0.0703809, -0.0832335, 0.0154163, -0.0057873, 0.0779768, -0.0236753, -0.0114421, -0.0476573, -0.0010590, 0.0136465, 0.0752500, -0.0443375, 0.0772168, 0.0081595, 0.1489798, 0.0991561, 0.0115904, 0.1983434, 0.0395799, -0.0184706, 0.1363550, 0.0031724, -0.0624186, 0.0399115, 0.0506258, 0.0287783, 0.0024279, -0.4808667, 0.0278093, -0.0732987, 0.0255355, 0.0270200, -0.0198608, 0.0312608, -0.2181814, 0.1118879, 0.0519991, 0.0178131, -0.0480703, -0.0265485, 0.1204475, 0.0974106, -0.0161309, 0.0279463, 0.0767297, 0.0221217, 0.0981063, 0.1145218, -0.0679343, 0.0197472, 0.2267244, 0.1638919, 0.0752007, 0.0197531, -0.0727337, -0.0080438, 0.0097427, 0.1420582, 0.1119991, -0.0958019, -0.0007137, 0.1099967, -0.0689616, 0.1077702, -0.0069677, -0.0241191, 0.0435674, -0.2705507, -0.2822470, 0.0752749, 0.1185725, 0.1685652, -0.4192066, 0.1634704, 0.4617664, 0.1965938, 0.1959372, -0.1774466, -0.0690006, 0.2033307, -0.0347321, 0.1531380, 0.2254974, -0.1815179, 0.2340192, 0.0981854, -0.2170269, 0.0361892, 0.0649950, 0.2626391, -0.1869117, 0.1769682, -0.1331562, 0.1602716, 0.3151225, 0.0318615, -0.0354331, -0.1715543, -0.3814526, 0.2272114, 0.1223313, -0.1781777, 0.2482991, -0.0410468, 0.3726221, 0.4882044, -0.1838085, 0.7125232, 0.4724791, -0.0140420, -0.0646924, 0.0219663, -0.5700171, -0.0306226, 0.3245635, 0.1604355, 0.2350401, -0.2641523, -0.1681978, 0.2031115, -0.1284361, 0.2199709, 0.1617279, -0.2816642, 0.2888219, 0.0884469, -0.3066518, -0.0191210, -0.0805698, 0.1779242, -0.2271637, 0.2587626, -0.0434045, 0.1818544, 0.2236807, 0.1909575, -0.0575309, -0.0976960, -0.5733433, 0.3270828, 0.2213064, -0.0670216, 0.1628148, -0.0199792, 0.4449277, 0.3866251, -0.2733011, 0.5557311, 0.3989047, -0.1744336, -0.1793787, -0.1514115, 0.0799666, 0.1048137, 0.2351380, -0.1073561, 0.0878576, -0.0046412, 0.0241350, -0.0632109, 0.0136065, -0.0921780, 0.0712459, -0.0621134, -0.1913496, -0.0383065, -0.1599261, -0.0261797, 0.2204176, 0.2214213, 0.0717768, -0.1217324, -0.0060639, 0.1272418, 0.1915897, 0.0257787, -0.1880144, -0.0895943, -0.0029749, -0.0730202, 0.0167039, -0.2073843, 0.1082940, 0.0007643, 0.0961888, 0.2238390, 0.0794077, 0.1598622, 0.2441006, 0.0851049, 0.2130300, -0.0580529, 0.0947029, 0.0127425, 0.0257957, -0.0596886, -0.1600253, 0.3398564, 0.1596936, -0.1375626, 0.0223206, -0.3097543, 0.0494726, 0.1904031, -0.0158551, -0.3471668, -0.3184298, -0.1933156, 0.0871454, 0.0619950, 0.1491055, -0.2577915, -0.0165791, -0.0320335, 0.2240953, 0.0840384, 0.0500197, 0.1428456, 0.1004140, -0.1867882, -0.1448863, -0.0774250, 0.1015324, -0.1198445, -0.1445405, 0.1829235, 0.0584519, -0.1814733, -0.0123247, -0.0365166, 0.0953681, -0.0426664, 0.0432775, 0.0085179, -0.0230134, -0.0765050, 0.0422760, 0.0564651, 0.1058885, -0.0566095, 0.1282128, -0.1125841, 0.0076965, -0.0020657, -0.0488287, -0.0887454, -0.0429257, -0.0508791, 0.1291589, 0.0175432, 0.0549796, -0.0862969, -0.0905309, 0.0244931, 0.0706463, -0.0519670, 0.0805046, 0.0415730, 0.0943323, -0.0629805, 0.0039024, 0.0317048, 0.0313667, 0.0383415, -0.1167270, 0.0057921, 0.0566920, -0.0372074, -0.0131852, 0.1564993, 0.1184280, -0.0518279, 0.0763402, 0.1259944, 0.0191402, 0.0065130, 0.0526330, -0.0916326, 0.0517125, 0.1163228, -0.0245695, 0.0324898, 0.0326282, -0.1219914, -0.0857200, 0.0983246, 0.0055346, 0.1284318, 0.0686674, 0.1399345, 0.0495971, -0.0225565, -0.1022654, 0.1238589, -0.1521411, -0.0785673, -0.0552174, -0.0839561, 0.0398359, 0.0149297, -0.1371358, 0.0208150, 0.1422793, -0.0087314, 0.0166419, 0.0322816, 0.0179972, 0.1156128, 0.0424566, 0.0636610, 0.1027110, -0.0846626, 0.1167852, -0.2298356, -0.2245020, -0.1123647, -0.0950886, 0.2066102, 0.2029307, -0.0170487, 0.2689619, -0.1633214, 0.1409250, 0.2149848, 0.2216823, -0.0433800, -0.1151589, -0.1841571, -0.0311754, 0.1093243, 0.1271717, -0.1219013, -0.1591097, -0.0447794, 0.0808155, 0.1908015, 0.0775067, 0.2417373, 0.1598247, -0.1139396, -0.0547357, -0.0147675, 0.1882911, 0.0083472, -0.2014997, 0.1608710, -0.1664989, -0.0689307, -0.2530954, -0.0526451, 0.1243577, 0.0504189, 0.0588898, 0.2409966, 0.1956516, 0.0655319, 0.1970404, -0.2232541, -0.0031053, 0.2110332, -0.1787072, 0.2251783, 0.0223252, -0.1602672, -0.1073640, 0.0744756, 0.0422986, 0.2562386, 0.0177157, 0.1085682, -0.0714417, 0.0609995, -0.0419816, 0.1714777, -0.0700824, -0.0793602, -0.1712700, -0.1937407, -0.0210907, 0.0743282, -0.0370424, 0.0339049, 0.1535102, -0.0307564, 0.1559739, 0.0745956, -0.0124169, 0.1940402, 0.1958417, 0.0066313, -0.0373003, -0.0471475, 0.0534952, -0.1287339, 0.0582062, -0.0470661, -0.4346946, 0.1242335, -0.1093059, -0.1703098, -0.0570967, -0.1964476, 0.0904282, 0.0260438, -0.0276017, -0.2490451, -0.1131799, -0.0746322, -0.0041550, 0.0780806, 0.1457092, -0.0823669, 0.0086352, -0.0367184, 0.1075761, -0.0264907, 0.0052090, 0.1032491, 0.0651261, -0.0092645, -0.0919687, -0.0497881, -0.0130053, -0.0710043, -0.0532862, 0.0902167, 0.0665948, -0.4005683, 0.1182049, -0.0435881, -0.0115679, 0.0160171, 0.0638931, 0.1050297, -0.0688651, 0.0408448, 0.0150345, 0.1057980, 0.0642475, 0.0746676, -0.0209498, 0.1485664, 0.0648646, 0.1804137, -0.0368001, 0.0440220, 0.1378322, 0.1742150, 0.0933884, 0.0667904, 0.0609428, 0.1149217, 0.1441496, 0.0202896, -0.0989071, 0.0164428, 0.0854039, 0.0891392, 0.1830612, 0.0707819, -0.1172743, 0.0558079, 0.0872285, 0.0476699, -0.0147259, -0.0922364, 0.0615690, -0.0468335, -0.1025803, 0.0173359, 0.1275039, 0.1927620, 0.3392452, 0.0446596, 0.4520833, 0.0248021, -0.1684541, 0.2647928, 0.1892020, 0.0396618, -0.0673803, 0.1361608, -0.2142612, 0.2364211, -0.2218919, 0.1890648, 0.2393332, -0.0014517, 0.4931085, -0.2398022, -0.0980378, -0.0834834, 0.0539522, 0.0552777, 0.4234270, 0.2087780, 0.1847177, 0.1111360, 0.3859698, 0.1300042, 0.1201611, -0.0888679, -0.1551738, 0.0734053, 0.2786045, -0.0157743, -0.0551540, -0.0477830, 0.3791983, -0.1381101, -0.0028975, 0.2964093, 0.3156513, 0.0593202, 0.2792980, -0.0155437, -0.0472798, 0.1558547, 0.2860335, -0.0154459, -0.0695142, 0.1530267, -0.1864331, 0.3264574, -0.2901360, 0.2390888, 0.1678359, -0.0352202, 0.3261464, -0.1404009, -0.0722414, -0.0809869, -0.0849118, 0.0167071, 0.3158000, 0.1295103, 0.2526712, 0.0085126, 0.2720937, 0.1919249, 0.0701646, -0.0655892, -0.1800836, -0.0859373, 0.1977984, -0.0099205, 0.0181188, -0.0440484, 0.3395770, 0.0378926, -0.0834524, 0.1728081, 0.2305374, 0.1709921, 0.3076050, 0.0368776, -0.1260579, 0.0613444, 0.1602380, 0.0592654, -0.0694327, -0.0520736, -0.1763894, 0.2110578, -0.2529200, 0.2072057, 0.0540198, 0.0843782, 0.3612466, -0.1582266, -0.0608436, -0.1841972, -0.0711978, 0.1378465, 0.1735812, -0.0664453, -0.0344291, -0.1382019, 0.2108558, -0.0244123, -0.0844510, -0.1620978, -0.0852388, -0.0728362, 0.1530182, 0.1137939, 0.0096506, 0.0227895, 0.3494776, -0.0066864, 0.1032873, -0.0324152, 0.1488666, -0.0287882, -0.0951775, -0.0666974, -0.0475533, 0.2321787, 0.2207931, -0.0086289, 0.1012503, 0.0623950, 0.0431161, 0.2919221, 0.1355352, -0.0088743, 0.0598625, -0.0100451, 0.0448614, 0.0954691, 0.1190778, -0.1041211, 0.1124418, -0.0153190, -0.0189279, 0.1921337, 0.0547959, 0.1523870, 0.1557945, -0.0426147, -0.1577599, -0.0166957, 0.1573036, 0.0025631, -0.1597901, 0.0468629, -0.0050053, -0.0995806, -0.2538108, -0.0499390, 0.1166713, 0.0596338, 0.1208092, 0.0136205, -0.0707211, 0.0132435, -0.1956115, 0.0424974, 0.1848064, 0.0981388, 0.1488691, -0.0671337, -0.0428495, 0.1831793, 0.1248239, 0.0743138, 0.0327251, 0.0201980, 0.0462715, -0.1084072, 0.0304272, -0.1815626, 0.0544362, -0.0387928, -0.1282624, -0.0443984, 0.0067757, 0.1898636, 0.1542090, -0.1458818, -0.1298359, -0.0509016, 0.1208363, -0.0182002, -0.1366182, -0.0694288, 0.0236075, -0.0146652, -0.0506069, -0.0256023, 0.1511094, 0.1974752, 0.3003988, 0.2247140, 0.1216212, 0.0704483, -0.0714591, 0.0511383, 0.1364945, 0.1507623, -0.2012311, 0.1149744, -0.2061449, 0.1372049, -0.2661009, 0.2872469, 0.1451021, 0.1219456, 0.3411378, -0.2426731, -0.2952712, -0.1288107, -0.1329077, 0.0568373, 0.0359931, -0.1521338, 0.1088114, -0.2086069, 0.2150555, 0.1532175, -0.1076525, -0.0179958, -0.0900751, -0.0997583, -0.0185211, -0.1385608, -0.0215105, 0.0576844, 0.1312060, -0.0074459, -0.1835173, -0.1002136, 0.0241855, -0.0972647, -0.2351202, -0.0895424, -0.0889154, 0.1339267, 0.1912087, 0.0942507, 0.2044731, -0.1600714, 0.1962833, 0.0583531, 0.1270717, -0.0844973, -0.1353013, -0.1078074, 0.0219059, 0.0628136, 0.0735329, -0.0879164, -0.0322407, 0.0391170, -0.0672954, -0.0143573, 0.0577081, 0.1495294, 0.0920501, -0.1180653, -0.1737313, -0.0136311, 0.1823887, 0.0718162, -0.2301812, 0.0571212, -0.0104378, 0.0617865, -0.2319501, 0.0036843, 0.1743676, 0.1949491, -0.0517503, 0.1179039, 0.4236422, 0.1806189, 0.0739904, -0.2263044, -0.1803805, -0.0089813, -0.3001890, 0.2469808, 0.0398473, -0.0635253, 0.0993451, 0.0474280, -0.1079261, -0.0095442, -0.0105596, 0.1242733, -0.3099894, 0.1748717, -0.1889786, -0.0086870, 0.3930613, 0.0563434, -0.2658998, -0.3230157, -0.2255361, 0.3257649, 0.2172606, -0.1538128, 0.0198776, -0.3111170, 0.4942210, 0.3306740, -0.1665065, 0.2573095, 0.4691561, -0.1679587, -0.4960174, -0.2107904, 0.1069121, -0.0341513, 0.0647925, -0.1401211, 0.1001067, 0.1391618, 0.1460237, 0.0118800, 0.0899839, -0.1413780, -0.0527263, 0.1761728, -0.0333811, -0.0404413, -0.2043808, -0.1279568, 0.0054710, 0.0986145, 0.0073583, -0.2254687, 0.0146063, 0.0733580, 0.0698618, 0.2392660, -0.0740920, 0.0565271, 0.0397667, -0.2161392, -0.1978439, -0.1663587, 0.1247211, 0.0232738, -0.0411697, 0.0486879, -0.0985735, -0.1735402, 0.1080784, -0.1558757, 0.1655712, 0.1782766, 0.0130647, 0.2326012, 0.0405238, 0.0897101, -0.1863036, 0.1577659, 0.0955603, 0.3138005, -0.1158005, 0.2562743, 0.0676404, 0.1667309, 0.0238127, 0.1451754, 0.0529260, 0.2480799, 0.2154320, -0.2319353, -0.2052281, -0.0725434, 0.2843393, 0.1161615, -0.2769919, -0.0604276, 0.1483517, 0.1249041, 0.0716608, 0.1821999, -0.1983997, -0.0834526, 0.2120049, 0.0922187, -0.0610261, -0.2032894, 0.0412954, 0.1751709, -0.0308019, -0.1676289, -0.0751029, -0.2918710, -0.0327703, -0.0945918, 0.2603569, -0.3893017, 0.3279219, 0.0577428, 0.0083571, -0.1342985, 0.0244298, 0.2729579, 0.0448048, -0.1043607, 0.0307805, -0.1239512, -0.0316290, -0.2511233, 0.1088148, 0.1395076, -0.1512850, 0.1291654, 0.2420044, 0.1523093, 0.2786264, 0.3584897, -0.1299082, -0.0174134, -0.1664097, 0.1747056, 0.2750815, -0.2541756, 0.2322697, 0.2700518, 0.2413839, 0.0349414, 0.1295878, 0.1484415, 0.2898600, -0.0735898, 0.1100143, -0.0888980, 0.2522220, -0.1466161, 0.0431653, -0.2526304, 0.0861837, 0.1015988, 0.2601342, -0.1439983, 0.0209178, -0.0000102, -0.1207696, 0.2435674, -0.1512321, 0.0296309, 0.0011871, -0.2678741, 0.1332975, 0.0792145, -0.0923030, -0.0570436, -0.2442441, -0.0797235, 0.1830003, 0.0888208, 0.1824234, -0.1385328, 0.1693616, 0.2313599, 0.0820394, -0.0750739, 0.0150910, -0.0034478, -0.1260551, -0.0242516, -0.1135563, 0.0601169, 0.0864055, 0.1453806, 0.0217231, -0.0046288, 0.1077608, -0.0419911, 0.4145041, -0.0693472, 0.1140103, -0.0091187, 0.0513359, -0.0891444, -0.0973827, 0.1898905, -0.0751561, -0.0042717, -0.0835169, 0.0924197, 0.0844486, -0.1175093, 0.1662159, 0.0422355, -0.1298343, 0.0027227, 0.0443418, 0.0154044, 0.3486033, 0.2570628, -0.1274582, -0.1802414, -0.0069632, 0.1463542, 0.2859408, -0.1611322, 0.0225201, 0.0304734, 0.3996117, 0.0637624, 0.0608305, 0.0417095, 0.4104267, -0.1711294, -0.1051114, 0.2392464, -0.0643548, 0.2127496, -0.2882258, 0.2276345, -0.0570898, 0.2612427, 0.1421988, 0.2389773, -0.0505243, 0.2027567, 0.2565438, -0.0291662, 0.2478877, -0.0632446, -0.0928351, 0.1403565, 0.3686572, -0.0980805, -0.1692412, 0.1243641, 0.3180739, 0.0330902, -0.2206016, -0.1701770, 0.2604132, 0.1576604, -0.0556080, 0.3173628, -0.3170278, -0.1982798, 0.3213958, 0.0207320, -0.2183691, -0.2021271, 0.2874293, 0.1551254, -0.3990541, 0.0459156, 0.1523553, 0.0990527, 0.0786802, 0.1375124, 0.0326073, 0.0720613, -0.2914521, 0.1463414, 0.1895981, 0.2264151, -0.0435813, 0.0011034, -0.0681324, 0.2046144, 0.0514937, 0.0010651, -0.0321771, 0.1201539, 0.1639055, -0.1541165, -0.0426513, -0.2261629, 0.1842456, 0.0201609, -0.1768213, 0.0349995, 0.0515869, 0.1468778, 0.1523486, -0.0395569, -0.2314358, -0.2202013, 0.1487015, -0.0254806, -0.0759235, -0.0989592, 0.0092130, 0.1530559, -0.0273558, -0.2477623, 0.0882095, 0.2336859, -0.0702076, 0.1728374, 0.2563248, 0.1218416, 0.0749192, 0.0082375, -0.1890032, -0.0748009, -0.3021032, 0.4171613, -0.0458153, 0.0221663, -0.0147499, 0.0374973, 0.0878286, 0.0265324, 0.0857672, 0.0349010, -0.1642538, 0.1396106, 0.1111680, -0.0046823, 0.2323572, 0.1814613, -0.0158852, -0.0593293, -0.1914144, 0.4021692, 0.2159274, -0.0820789, 0.0055811, -0.1004677, 0.2186196, 0.0106773, 0.1736907, 0.1413342, 0.2177635, -0.1681282, -0.3718553, -0.0038361, 0.0739158, 0.0566773, -0.1393455, 0.0718275, -0.0070234, 0.0254869, 0.0472016, 0.0912500, 0.0914199, -0.0765151, 0.0658635, 0.0727319, 0.0277393, 0.0040502, -0.0097737, 0.0248489, -0.0507617, 0.0406708, 0.1091295, -0.0179237, -0.0301415, 0.0330453, -0.0566480, -0.0886815, -0.0297173, 0.0648158, 0.0832814, -0.0621271, -0.1680482, 0.0434127, 0.0448304, -0.0191164, -0.0847299, 0.0549264, 0.0015091, -0.0020976, -0.1221277, 0.0613076, 0.0827847, 0.0547523, -0.0224335, -0.1099267, 0.1211955, 0.1132369, 0.0698487, 0.0076269, -0.1712370, -0.1413330, 0.0939804, 0.0069555, 0.1387924, -0.0775671, 0.1871460, 0.0031111, 0.0195456, -0.0421972, 0.0144851, 0.0612710, 0.1843702, 0.2377636, 0.0224646, 0.0769347, 0.1880356, 0.0503082, 0.0110602, 0.0410768, -0.0665435, 0.0796013, 0.2348715, 0.2312932, -0.1947388, 0.0484256, 0.1999324, 0.2480163, 0.0796974, -0.0218422, 0.1181810, 0.1090780, -0.1567667, -0.0104600, 0.0820444, 0.1352636, 0.0917321, -0.0919191, 0.0155196, 0.1850895, 0.3566609, 0.2155797, -0.0638111, 0.1908010, 0.0051207, 0.1160108, -0.0019641, 0.0080649, -0.1013552, 0.0552870, 0.3091822, -0.0938511, -0.2107424, -0.2182567, 0.2411147, 0.0103776, -0.1507278, 0.1319754, 0.2250119, -0.0223088, 0.0386480, 0.2122533, -0.2460057, -0.4739778, 0.3599423, 0.1536336, -0.1135438, -0.1831983, 0.0284197, 0.2412601, 0.0074522, -0.2193597, 0.3136828, 0.2173650, -0.1147258, 0.2264964, -0.0274465, 0.1985195, -0.0915011, 0.1998129, -0.0198498, 0.2502999, -0.0218470, 0.0329525, 0.2107139, -0.1863336, 0.1932705, 0.0864200, -0.0826152, 0.2095272, 0.3147561, -0.0846316, -0.1177840, 0.0839876, 0.2314124, 0.1552679, -0.1292303, -0.1787980, 0.0714750, 0.0982051, -0.0965609, 0.1043090, -0.1181459, -0.0878221, 0.1062246, 0.0412072, 0.0120703, 0.1797840, 0.1514922, 0.1935493, 0.0935457, 0.0081697, 0.0360622, -0.2692896, -0.2800792, -0.2275594, 0.1691001, -0.2253736, 0.3374147, -0.0852970, 0.1171736, -0.0865330, 0.2244384, 0.1678799, -0.0139080, -0.0120317, -0.1174496, 0.0408868, -0.2837943, -0.3409690, 0.2834657, 0.1377059, -0.1386566, -0.0513742, 0.0662854, 0.1458604, 0.2363875, 0.1319511, -0.0501631, -0.1720477, -0.1972721, 0.1383830, 0.1389266, -0.3308575, 0.3252095, 0.3215220, 0.0282892, 0.0402558, 0.1029100, 0.1826589, 0.1354731, 0.0992420, 0.3106563, -0.2098039, 0.0931489, -0.2201869, 0.0022471, -0.2760627, 0.2722426, -0.1163729, 0.2411959, -0.0274136, 0.1832406, -0.0502269, -0.1729994, 0.1637068, -0.2166429, 0.1638324, -0.1120639, -0.3389325, 0.0938779, 0.1840971, -0.1289443, -0.1995082, -0.1465880, 0.0913730, 0.0524281, 0.0575521, -0.1505949, -0.2071012, 0.0362177, -0.0730642, -0.0001249, -0.1674736, 0.3574713, 0.1936473, -0.1542685, -0.0554032, -0.0207822, 0.2063252, 0.0287339, 0.1599535, 0.2276932, -0.0992537, -0.1826025, -0.1496420, 0.2973740, -0.0221892, 0.1695059, -0.1129001, -0.2746725, -0.0453669, -0.0179990, 0.1993562, -0.0368067, -0.1221195, 0.1635991, -0.0076058, -0.1005548, -0.1621026, -0.1282490, 0.1731222, -0.1756081, 0.0943469, 0.0564398, 0.1776090, 0.2219814, 0.3716842, -0.4603519, -0.0850742, -0.2703945, -0.0084275, 0.2882864, -0.2355915, 0.0324463, 0.1141126, 0.4410161, 0.3195011, -0.3111375, 0.2550853, 0.2300459, -0.3711510, -0.0937150, 0.4208469, 0.0336900, 0.3076217, -0.2463459, 0.5553921, -0.0412793, 0.2089218, -0.1752362, 0.2429176, -0.0909241, 0.3008813, 0.4540476, -0.1196509, 0.5136747, 0.1163765, 0.0899673, 0.3435031, 0.1843425, 0.0160951, -0.0674560, 0.2535917, 0.3168913, 0.0737301, -0.2131352, -0.0640465, 0.2049358, 0.2212691, 0.0646861, 0.2644549, -0.0965548, -0.0075308, 0.2671807, -0.0461153, 0.0264967, -0.0554884, 0.1762841, 0.2056948, -0.3305044, -0.0025188, -0.0804488, 0.0866264, -0.0158886, 0.0880453, 0.0166706, 0.1209548, -0.1557277, 0.0752222, -0.0186569, 0.1406814, -0.0724294, -0.1202993, -0.0120846, -0.0469668, -0.0805431, 0.0513948, -0.0543704, 0.1120353, 0.1169628, -0.0668628, -0.0113028, -0.0827445, 0.0719676, 0.1319835, -0.1124472, -0.1319417, -0.0325448, 0.0228730, 0.0376107, -0.1240707, -0.2193330, -0.0772852, 0.0115943, -0.0562809, 0.0020916, 0.0495954, 0.0354306, 0.0859134, 0.0372484, -0.0198672, 0.0301407, 0.4749477, 0.0659718, 0.3493434, 0.1338158, 0.4322615, -0.1990350, 0.2172019, -0.0673993, 0.2566860, -0.2741736, 0.0422815, 0.0898568, 0.0123280, 0.1022025, -0.0101340, -0.0707715, 0.3146263, 0.3280056, -0.0180060, -0.0697337, -0.0091047, 0.1471724, -0.0269007, -0.0498981, -0.1623898, 0.2090189, 0.1514826, 0.1551129, 0.1399688, -0.2075785, -0.1098598, 0.0771334, -0.3124045, 0.0540717, 0.1815807, 0.1797170, 0.2539734, 0.2604646, -0.1986277, -0.3202823, -0.1222381, 0.0778499, 0.0635034, -0.0396658, 0.0647980, -0.0378017, -0.0012209, 0.0032619, 0.0426529, 0.0355147, -0.0327521, 0.1025354, 0.0152277, 0.0305709, -0.0039325, 0.0133206, 0.0529063, -0.1545769, 0.0924239, 0.0544394, -0.0008190, -0.0409146, -0.0031173, -0.0136198, -0.0056963, -0.1613562, 0.0269650, 0.0570627, -0.1080438, -0.1221460, 0.0331622, 0.0913213, -0.0836853, -0.0166034, 0.0669564, -0.0291652, 0.0330487, -0.0427389, -0.0073994, 0.0543740, 0.0416817, 0.0579177, -0.0839381, -0.0537580, 0.1088500, 0.1195515, -0.0441509, -0.1040339, -0.1288288, 0.1341710, 0.0143798, 0.1094862, -0.0610564, 0.0767439, 0.0489499, 0.1120636, 0.0419022, -0.1805692, 0.1406534, 0.3834932, 0.1676146, 0.0264064, -0.0054104, 0.1089106, 0.0505508, -0.0877325, 0.1791348, 0.0471935, 0.0011543, 0.2646769, 0.2202672, -0.1113584, 0.0350782, 0.0962337, 0.1219548, 0.0248214, -0.1964010, -0.0236494, 0.1006940, 0.0096465, 0.3662162, -0.0145768, 0.4125103, 0.1227103, 0.4007570, -0.1393981, 0.2458024, -0.0532448, 0.3109244, -0.2706940, 0.2379119, 0.2930983, -0.0876713, 0.0872493, -0.0517661, -0.1322842, 0.3582015, 0.4258492, -0.1855724, -0.2660764, -0.0193489, 0.1912157, 0.0572479, -0.3013873, -0.2299276, 0.1770097, 0.0283545, 0.0717552, 0.3050174, -0.3234530, -0.3447818, 0.2908188, -0.1813868, 0.0383754, -0.1715488, 0.1875895, 0.2722600, -0.0058759, -0.2316539, -0.0102389, 0.1805601, 0.0097890, 0.1342532, 0.0200923, 0.1098894, -0.0263365, -0.0836959, 0.0952206, 0.2554839, -0.0513132, 0.0466313, 0.0814923, -0.0563207, 0.1599315, 0.1539235, -0.0789307, 0.0915855, 0.0865477, -0.1104073, -0.2378905, 0.0092620, 0.0608132, 0.2031681, -0.3080954, -0.2601213, 0.0736910, -0.0314080, 0.0519070, -0.0520482, -0.1484409, -0.0785666, 0.0889827, 0.0796754, 0.0351804, -0.0288576, -0.1111901, 0.2874953, 0.1549047, -0.0511936, 0.0127074, 0.1825616, 0.0089556, 0.2241292, 0.2573323, 0.1292355, -0.1984332, 0.1986365, 0.0715502, 0.2016957, -0.0613882, 0.1091896, -0.0853100, 0.1057813, -0.0163673, -0.0177234, -0.0378278, 0.1904945, 0.3692907, -0.2426842, -0.1264121, -0.1168695, 0.3138804, 0.1621710, 0.1725549, 0.0250663, -0.0005135, 0.1113268, -0.0055379, -0.0166504, 0.0553821, -0.2155102, 0.0908080, 0.1109132, 0.2096964, 0.0552251, 0.1066875, 0.1727903, 0.2407918, -0.2147188, 0.0435150, -0.0736497, -0.0913212, -0.0997085, -0.0184951, -0.0653589, 0.1960386, -0.0231378, 0.2425284, 0.3031689, 0.3680361, 0.0778798, -0.1045645, -0.1047851, 0.0696028, 0.2970327, 0.0680506, 0.0004003, 0.4205916, -0.0638179, -0.0180961, 0.0489463, 0.0247970, 0.4550981, 0.0237524, 0.0019698, 0.1471620, 0.0398601, -0.0331605, -0.0667370, -0.0237013, -0.1030572, 0.2738847, 0.2944533, -0.0716346, -0.0481973, -0.1607058, 0.2749546, 0.0000204, 0.1613192, 0.3001739, -0.2006657, 0.0466810, -0.0639341, 0.3228562, -0.1070002, 0.0005073, 0.2754988, -0.0990788, -0.0857161, 0.0619063, 0.0887170, -0.0142222, 0.2550688, -0.0436781, -0.0014800, 0.0868122, -0.0898105, 0.1079178, 0.1844196, 0.1429679, -0.0775897, 0.2625698, 0.2069211, 0.5472116, 0.5328961, -0.1985298, 0.1734169, 0.0330683, 0.1133092, 0.2557769, -0.2552532, -0.0386182, 0.1765600, 0.4726398, 0.2793897, -0.0882327, -0.0331910, 0.3022054, -0.3407491, 0.1116923, 0.1691501, 0.0394966, 0.0826047, -0.0770265, 0.2495084, 0.0387738, -0.0254990, -0.0991439, 0.2393852, -0.0837346, 0.4412478, 0.2949217, -0.0322172, 0.4099075, -0.0087281, 0.0916740, 0.3551217, -0.0953003, 0.0099942, -0.0761509, 0.2517877, 0.4120229, -0.0282274, -0.1582441, 0.2226274, 0.1064334, 0.1493686, -0.0031331, 0.2809645, 0.1895067, 0.0201457, 0.1764870, 0.0985613, 0.1796486, -0.1026363, -0.1089974, 0.1114570, 0.0168537, -0.3823063, -0.2844009, 0.0051018, 0.0120268, 0.0560601, 0.1034791, -0.0095557, -0.0917645, -0.1606146, 0.0112651, 0.1478595, -0.0822327, 0.0186515, -0.1240488, 0.0921716, -0.0870091, 0.1256172, 0.0619088, 0.0752378, -0.0178935, 0.0017987, 0.0185457, -0.0546096, 0.0561888, 0.1147712, -0.0972393, -0.0101994, -0.0991243, -0.0319741, 0.1048044, -0.2040623, -0.1714600, 0.0416429, -0.0211343, -0.0174092, 0.0993737, -0.0187731, -0.0207297, 0.0465188, 0.1515521, -0.0624829, -0.0442505, 0.1806968, 0.0389140, 0.2113922, 0.1101748, 0.1322725, -0.0388672, 0.0744510, -0.0311853, 0.1953299, -0.3154835, 0.1465063, 0.0718917, 0.0383081, 0.0911085, 0.0596817, -0.0017177, 0.2257629, 0.1178272, -0.0359246, -0.2376652, -0.0126618, 0.0410707, -0.0782316, -0.0511099, 0.1174139, 0.0772996, -0.0240775, 0.0117524, 0.0646584, -0.0738400, -0.1084998, 0.1264487, -0.2296365, 0.1350838, 0.0036149, 0.0664540, 0.1775237, 0.1423277, -0.1941302, -0.2809217, -0.0351576, 0.0397719, 0.0160374, -0.0828539, -0.0013842, -0.0625366, -0.0758253, 0.0904641, 0.1395570, 0.0883799, 0.0887538, 0.0252070, 0.0921814, 0.0488668, 0.1602068, 0.0573310, 0.0762435, -0.1149362, 0.0111880, -0.0711996, -0.0008560, -0.0188056, 0.1045406, -0.1632361, 0.0580689, -0.0246393, -0.0479392, 0.0466178, -0.1177751, -0.1671406, -0.0500292, 0.0782095, -0.0007973, 0.0365532, -0.0272369, -0.1164222, 0.0900290, -0.0907879, -0.0328303, 0.0145110, -0.0581686, 0.0529393, -0.1701630, 0.0054158, 0.0062154, 0.1463661, -0.1053535, -0.0127070, -0.0076949, 0.1446386, 0.0614416, 0.0201816, 0.0377510, 0.1731476, 0.1312188, 0.1120735, -0.0477243, -0.3190657, 0.1727637, 0.1504233, 0.1357550, -0.0030060, 0.0348121, 0.0266117, 0.2204321, -0.2015669, 0.0685930, 0.0211281, -0.1840223, 0.1956341, 0.1191981, -0.0737235, 0.1265120, 0.1824350, 0.0450891, -0.0754176, -0.0532362, -0.0230069, 0.0473874, -0.0503188, 0.1854431, -0.0468569, 0.2834034, 0.0507697, 0.3134167, -0.1033919, 0.1758690, -0.1115806, 0.1849289, -0.3006316, 0.3827335, 0.3738714, 0.1704911, 0.3834264, -0.0257199, -0.0768981, 0.2910868, 0.1601702, 0.0306511, -0.2549221, 0.0540083, 0.3519988, -0.0321617, -0.2413903, 0.1576842, 0.1499328, 0.1241573, -0.0363129, 0.2623649, -0.0754890, -0.2034402, 0.3430054, -0.1638152, 0.1069963, -0.0672225, -0.0268526, 0.3337823, 0.0842881, -0.5477886, -0.3410802, -0.0780127, 0.0064252, -0.0489638, -0.0849749, 0.0184488, 0.0821086, -0.0764014, 0.0293961, -0.0410667, 0.0406332, 0.0164982, -0.0238394, 0.0009182, -0.0308937, -0.1346903, -0.0800997, -0.0772550, 0.0455907, 0.0558563, -0.0694579, 0.0511294, 0.0351096, -0.0979499, 0.0313577, -0.0246664, 0.0560355, -0.0208149, -0.0761011, 0.0376486, 0.0444432, -0.0120413, 0.0386983, -0.0464265, -0.0036856, -0.0262326, -0.0057702, 0.0410555, -0.0288182, -0.0161921, 0.0048418, 0.0242448, -0.1249447, 0.1600865, 0.1229583, 0.0902464, 0.0876502, 0.0831791, 0.0434269, 0.0644763, 0.2229599, -0.1624908, -0.0322852, -0.1864532, -0.0394388, 0.0398137, -0.1021349, 0.1144634, 0.1888604, 0.0484390, 0.0920126, 0.2119238, 0.1216233, 0.1850482, 0.1367357, -0.0781609, 0.0285710, 0.1701656, -0.0648396, 0.0246426, 0.0708206, -0.0079330, 0.1580162, 0.0615315, 0.0498609, 0.1060068, 0.0511675, 0.1838958, 0.1640264, 0.2869260, 0.1105984, 0.3953545, 0.0996647, 0.2165896, -0.2048649, 0.4663979, -0.1046685, 0.4401844, -0.1199366, 0.0455386, 0.1143474, 0.1512172, 0.3061185, -0.0431636, 0.1567135, -0.1926660, 0.1362356, 0.1869920, 0.5371080, -0.0307674, 0.2584867, 0.5059863, 0.0779352, -0.1471652, 0.1206644, -0.1309894, 0.3569628, 0.4127564, 0.0741535, 0.4578399, 0.2019666, 0.2356907, -0.0153862, -0.2404052, -0.0312343, 0.0190977, 0.3815177, 0.0892154, -0.0545236, 0.1296338, -0.1686929, 0.1017634, 0.0682292, -0.2126291, -0.0164304, 0.1485715, -0.1826223, 0.4704595, 0.1517623, -0.2356967, 0.6250950, -0.2250502, 0.0727888, 0.0644388, 0.1137609, -0.1158936, -0.0380627, -0.1877245, 0.2674817, 0.0656524, 0.4832686, -0.0600204, 0.0509768, 0.0021504, 0.5189722, 0.2395429, 0.0957364, 0.7467171, 0.0858230, 0.0672635, 0.2827207, 0.1204741, -0.1650231, 0.0595181, -0.0585302, 0.4046339, 0.0966766, -0.2124218, 0.0126055, 0.0721681, 0.1412120, 0.0679560, 0.0177551, -0.1038687, 0.2270511, 0.0596723, -0.0084831, 0.1240769, 0.1135985, -0.0946607, 0.0574974, 0.0500736, 0.2112502, 0.0778415, 0.3599213, -0.0825495, -0.1862487, -0.0303958, -0.0446935, 0.1433026, -0.0050898, 0.0695975, 0.1411228, 0.0455728, 0.2141601, 0.4179088, 0.0553032, 0.1093840, 0.0215256, 0.0881670, 0.2487791, -0.1374958, 0.1339301, 0.1216539, 0.1977522, 0.2189902, -0.1775504, 0.1693432, 0.1978890, -0.1916279, 0.0141557, 0.0348659, -0.0510607, -0.3336484, 0.2547331, -0.0927851, 0.1004287, 0.1421144, 0.0047033, -0.2482178, 0.2198757, -0.0220641, 0.0310028, -0.0061982, -0.0394243, -0.2521432, -0.1958906, -0.3715267, 0.2081291, 0.0298488, 0.0425015, 0.0136313, 0.0445131, -0.0146048, 0.5134400, 0.1131417, 0.0889454, 0.1306831, -0.1363013, 0.1533057, 0.3831161, -0.1260949, -0.0093756, 0.0911617, 0.0479725, 0.4187593, -0.0026269, 0.1213451, 0.3099106, -0.0344873, 0.0504321, -0.1389172, 0.2105670, 0.1875823, 0.0558545, -0.1538961, 0.1185253, -0.2659825, 0.0343474, 0.1148340, -0.1784109, 0.1685192, 0.0892871, -0.0788431, -0.1384851, 0.1145356, 0.1270817, 0.1174032, -0.0373600, 0.1820998, -0.0366519, 0.0602864, -0.1325451, -0.0046881, -0.2641541, -0.0978234, -0.0741055, -0.3210647, 0.1834671, 0.0094369, -0.1323747, -0.0082675, 0.2090026, -0.0828090, 0.0257060, -0.0317095, -0.0404640, 0.1331793, 0.0680630, 0.0342875, 0.0539565, -0.1121321, 0.0463647, -0.1020501, 0.0422331, -0.1670570, 0.0539880, -0.0771540, 0.0544261, -0.0295544, 0.1256784, -0.1211872, -0.0771928, -0.0364397, -0.1618955, 0.0107047, -0.1410439, -0.2187970, 0.0931879, 0.1000323, -0.1779136, -0.0816540, -0.0963412, -0.0041639, 0.1410743, -0.1304673, -0.0976894, -0.1667281, -0.0553557, -0.1513846, 0.0288983, -0.1366629, 0.1031370, -0.0198495, -0.0568440, 0.0766725, -0.0655885, 0.0728781, 0.0653046, 0.0017099, 0.0957227, -0.1935588, -0.0843454, -0.0099259, 0.1084491, -0.1056303, 0.1566460, -0.2141992, 0.2010716, 0.1052062, 0.1476163, -0.0020039, -0.1017982, -0.2531111, -0.1736681, 0.1941820, 0.0291971, -0.0611425, 0.1511690, 0.0399089, 0.0053218, -0.0544371, 0.0409578, 0.2505790, 0.0297524, 0.0472983, -0.0170941, -0.1861376, -0.1207490, -0.0472189, 0.0946949, -0.1309268, 0.1850135, 0.2375684, 0.1041454, -0.0102710, 0.0218701, 0.1518147, 0.1248695, 0.1652853, 0.2782801, -0.0638805, 0.1046317, 0.0495651, 0.0023592, 0.0185070, 0.0880485, -0.0474914, 0.0003702, -0.0861405, -0.1304790, 0.1899589, 0.1111229, -0.0069156, 0.1262878, -0.0525736, 0.0794487, 0.1129845, -0.2321674, 0.1708546, -0.0313479, 0.1863007, 0.0626795, -0.0432257, -0.0194243, 0.1409807, -0.0830909, 0.0138531, 0.0330894, 0.0184050, 0.0636402, 0.0187219, 0.1204299, -0.0020146, 0.1202533, -0.0063634, -0.0340639, -0.0231065, -0.0160524, -0.0956124, -0.0712608, 0.0979203, 0.0508607, -0.0218548, -0.0360614, 0.1105435, 0.0214932, 0.0826901, -0.1868355, -0.1923797, 0.0999359, -0.0662290, 0.1527715, -0.1116618, 0.1214289, -0.3289790, -0.0440600, -0.0847223, 0.0723310, 0.1170337, 0.0715863, 0.0258351, -0.0485325, -0.1342838, 0.1560736, -0.0739471, 0.1202931, 0.1010130, -0.0004979, 0.1013047, 0.1729119, 0.0430695, -0.1448455, -0.0446967, -0.1006525, 0.1234420, 0.1482229, -0.0347221, -0.0225141, 0.0718165, -0.0132606, 0.1170482, 0.2120907, -0.0296344, -0.0029151, 0.0655058, -0.0586040, 0.0835240, 0.1909943, 0.1096300, 0.1778256, -0.2112495, -0.0276342, 0.2638637, 0.0159200, 0.2099580, -0.1559254, -0.0584402, 0.1875303, 0.0914082, 0.0619179, -0.0688975, -0.4207382, 0.0317818, 0.1081795, -0.0771821, 0.2807870, -0.0253223, 0.2646498, -0.0293104, -0.0812056, 0.0504589, 0.0208236, -0.0819665, 0.0412808, 0.3280714, -0.0341781, 0.2564686, 0.1073847, 0.1640624, 0.0390962, 0.3114112, 0.0056216, 0.1416835, -0.1329249, 0.2625118, 0.0317535, 0.3520522, -0.0160278, 0.0693117, -0.0118555, 0.1049574, 0.2544609, -0.1042073, 0.2511132, -0.0652732, -0.1558304, -0.0168469, 0.6371496, 0.1189664, -0.0281543, 0.3404281, -0.1863487, -0.1917165, 0.1253169, -0.3063981, 0.5209503, 0.1892276, 0.0308751, 0.4538743, -0.0464464, 0.1348474, 0.1676605, -0.2218577, -0.2544844, 0.0916446, 0.2590738, 0.2729964, 0.0369147, 0.2449245, -0.0537089, 0.0105736, 0.0629244, -0.1192439, 0.0112393, -0.0116049, -0.1958085, 0.2928809, 0.0909461, 0.0425542, 0.0559263, -0.2907033, 0.0089675, 0.1697677, 0.1061079, -0.0648398, -0.3646671, -0.2673969, 0.2413063, 0.0633880, -0.0467134, -0.3642220, -0.1061376, -0.0441495, 0.1506564, 0.1073753, 0.2180953, 0.1003773, 0.0377370, -0.0648685, -0.0904552, -0.1962233, 0.1537526, -0.0872988, -0.1695780, 0.2386219, -0.0416102, 0.0895398, 0.0580457, -0.0682681, 0.1387184, 0.0474926, 0.0714240, -0.0505276, 0.0919497, 0.0159677, -0.0401286, 0.0296550, 0.0565681, 0.0469560, -0.0228224, 0.0784439, 0.2651875, 0.0516308, 0.0761399, -0.1304941, -0.0429466, -0.0287128, 0.0630951, 0.1233458, -0.0388977, -0.0363487, 0.0329443, -0.0687603, 0.1424897, 0.1419525, 0.1098688, 0.0036196, -0.0394596, 0.0664709, 0.0512434, -0.0860952, 0.0652121, -0.0728112, 0.0195103, 0.0383249, 0.0058243, 0.0915653, 0.0424149, -0.0062912, 0.0818615, 0.0883557, -0.0907699, -0.4450717, 0.1431894, 0.0326986, -0.1947941, 0.3799845, -0.0042310, -0.1134195, 0.4295031, -0.3302402, 0.0297977, 0.0691920, 0.0720063, -0.2767107, -0.2982760, -0.3505269, 0.2785596, -0.0250866, 0.1851568, -0.1137144, -0.0384673, 0.0127281, 0.4061829, 0.0709890, 0.1511977, 0.3860765, -0.0492099, 0.0008588, 0.2010982, -0.0833669, -0.1574974, 0.0230554, -0.0947336, 0.4082361, 0.0305731, 0.0020838, 0.1570048, 0.0531874, 0.0827143, -0.2542651, 0.0529389, 0.1594259, 0.0617528, -0.0890670, 0.1822296, -0.1793151, 0.0517113, 0.1925389, -0.0348087, 0.0810427, 0.1730097, -0.2622335, -0.0419288, 0.0223861, -0.0480091, 0.1083340, -0.0344944, 0.2573018, -0.0729829, 0.0357387, -0.1094531, 0.1202139, -0.1276901, -0.0819583, -0.1853430, -0.1708098, -0.0396315, 0.0011097, -0.1643048, -0.0433540, 0.3267112, 0.0111268, -0.0232869, 0.0877330, 0.0325565, 0.2090624, 0.0887489, 0.0778469, 0.1788665, -0.0274480, -0.0810517, -0.1925074, 0.0545654, 0.0417672, -0.0983626, 0.0918253, 0.0281199, 0.0100439, 0.1857399, -0.3572949, 0.1276060, 0.1087161, 0.2333337, -0.1160005, -0.3033823, -0.1406098, -0.0367976, 0.0279704, 0.0641951, -0.2072954, 0.0208076, 0.0564245, 0.2052140, -0.0500717, -0.1061150, 0.0864435, -0.0043929, -0.1863321, -0.0760081, -0.1016538, 0.0074291, 0.0042162, -0.0232747, 0.4055842, -0.1354635, 0.0837575, 0.1188467, -0.0555713, 0.0436675, -0.2616045, -0.0065227, 0.1122476, 0.1793838, -0.1720557, 0.3190882, -0.2128503, 0.0843781, 0.0611383, 0.0404127, -0.0028935, -0.0450712, -0.1044599, -0.3594344, 0.0237148, 0.0217792, 0.0433454, -0.0412878, 0.1946539, 0.0333381, -0.0551442, 0.0580220, 0.2171507, 0.0220341, -0.0023251, -0.3947675, -0.2001158, -0.0875233, -0.0707203, 0.0027920, -0.1091397, 0.2610102, 0.1816382, 0.1606393, 0.1110787, 0.0781281, 0.0790229, 0.2356168, 0.0979780, 0.1854203, -0.0776648, 0.0721352, 0.0113695, -0.0840642, 0.0193635, 0.0898691, -0.0106550, -0.1059722, -0.1226372, -0.0372523, 0.1641017, 0.2970653, -0.1316246, 0.0626846, -0.0571872, 0.0447470, 0.0254956, -0.0956633, 0.1407951, -0.0061936, 0.2706836, 0.0917491, -0.1580313, 0.0131169, 0.0296879, 0.0564182, 0.0046555, -0.0172873, 0.1511331, 0.0842964, 0.0325762, 0.0712602, -0.0462619, 0.0619232, -0.0120956, 0.0436336, -0.0037761, -0.0781409, -0.0088394, -0.0258696, 0.2750287, -0.0137274, -0.1069729, -0.0119406, 0.1627479, -0.2127193, 0.4045681, -0.0732816, -0.1569914, 0.3223040, -0.1742705, 0.2076454, 0.1029467, 0.2418482, -0.3431051, -0.2401314, -0.2068824, 0.3547107, 0.0133602, 0.2548304, 0.0320556, -0.0944727, -0.0724398, 0.3389701, -0.1412135, 0.2774028, 0.4852117, 0.0214332, 0.2078706, 0.2302893, 0.0683486, -0.0914367, -0.0721417, -0.1376995, 0.3949804, 0.1771103, 0.0398217, -0.0344554, 0.1816011, -0.0439427, 0.0004442, 0.2093097, 0.0166809, -0.0376381, 0.0048508, -0.0361368, 0.1361021, 0.2857335, 0.1864360, 0.1495298, -0.2714364, 0.1413390, 0.2082880, 0.0555956, 0.1469997, -0.1680798, -0.0411878, 0.2819906, 0.1719893, 0.0496993, -0.1493427, -0.2867637, 0.1012429, 0.0364864, -0.0062393, 0.0053512, -0.0421151, 0.2936685, -0.1889739, -0.2701332, -0.1084913, 0.2331343, 0.0158004, -0.1083285, 0.2214420, -0.0725741, 0.2396041, 0.0452047, 0.1813311, 0.2691153, 0.0144177, 0.0796965, 0.0234621, 0.0379822, -0.0187648, 0.1584746, -0.2394365, 0.2506056, 0.2420950, 0.0755866, -0.1419590, 0.0109313, -0.1390290, -0.1764102, 0.2544899, -0.0946356, -0.0613822, 0.3633536, 0.1128559, -0.0800020, -0.0096516, -0.5064907, 0.1021852, 0.0134526, -0.1736181, 0.3070951, -0.3587470, 0.0231053, 0.0688493, -0.1675603, -0.0361254, 0.1677283, 0.0181391, -0.0713002, 0.1359941, -0.0641336, 0.4956893, 0.0755435, 0.3179151, 0.1136985, 0.0025147, 0.0065452, -0.1321746, -0.1522667, 0.0007875, 0.0105971, 0.1434909, 0.1707175, 0.0120716, 0.1065346, -0.1455475, 0.1597212, 0.1200386, 0.1346045, -0.0082952, -0.2203089, -0.1565679, 0.2312870, 0.0890816, -0.0402669, -0.0875556, -0.0576493, -0.0818980, 0.0310465, -0.0383581, 0.1043909, 0.0111909, 0.0906653, 0.0033753, -0.0762641, -0.1597565, 0.2473729, -0.0180029, -0.2004188, 0.0376851, -0.0318235, 0.1055412, -0.1002424, 0.0866864, 0.1254513, -0.0861105, 0.1052199, 0.1082567, 0.0892045, -0.0447438, 0.1454587, -0.0116248, -0.1890116, -0.0388580, -0.1256440, 0.1980920, 0.5996550, -0.1986762, -0.1154632, -0.3371731, 0.0784509, 0.0597334, 0.0096606, 0.2202944, 0.0698231, 0.3090981, 0.0024781, -0.3761886, 0.0233109, -0.0807571, -0.0027341, -0.0849626, 0.0803651, 0.3193519, -0.0129889, 0.0542720, 0.2191400, -0.2328994, -0.0338800, -0.0060959, 0.2149777, 0.0649841, 0.0833286, 0.1144091, 0.1278524, 0.0868385, 0.0713293, -0.0595325, 0.2150695, -0.0585626, -0.3717602, 0.4493287, -0.0310164, -0.1248037, 0.2257132, -0.3782470, 0.0262357, 0.2208528, -0.0306312, -0.3043706, -0.2188894, -0.1997776, 0.3023874, -0.0203697, 0.2770370, -0.1614403, 0.0310374, 0.0082725, 0.3041136, 0.0592840, 0.1361492, 0.4569908, 0.1265771, -0.1432994, 0.1149376, -0.0543883, -0.1377264, -0.0198754, -0.0201399, 0.2780262, 0.1962465, -0.3513069, 0.2131081, 0.0338645, 0.1100909, 0.0497124, 0.0894244, -0.0138472, 0.1119117, -0.0151253, -0.0569929, 0.1966311, 0.1803258, 0.0711852, 0.0728792, -0.1050462, -0.0953577, 0.1355404, -0.2611713, 0.0405403, -0.0642892, -0.1245473, 0.3637606, -0.2288057, -0.1101901, -0.1421526, -0.1549436, 0.0630290, 0.2260325, -0.1573795, 0.1113998, -0.0652892, 0.0984886, 0.1216200, -0.0431790, -0.0389725, -0.0805000, -0.0013188, -0.0580885, 0.1315262, 0.0119873, 0.0680910, 0.1967815, 0.1947466, 0.1120369, 0.1162162, 0.0390531, -0.1913650, 0.1497918, 0.1227660, -0.2428756, 0.2207988, 0.0082404, -0.0857152, 0.2789183, -0.2178800, 0.0220586, 0.1930984, 0.2175172, -0.0358245, -0.0376138, -0.0971791, 0.1009399, -0.0574463, 0.1338677, -0.1545877, 0.0827546, -0.0147762, 0.2194646, 0.1052716, 0.0677795, 0.3377716, 0.0779485, -0.0843323, 0.2523557, -0.0029902, -0.1152820, 0.0272761, 0.0988264, 0.2208458, -0.0616275, -0.1059828, 0.0628307, -0.1321607, 0.0465654, 0.1575500, 0.1381961, 0.1552071, 0.2420451, 0.0328161, -0.2597761, 0.2173453, 0.0423094, -0.0258847, 0.0146357, -0.2377851, -0.0974717, 0.0774199, -0.3370609, -0.0247404, -0.1418457, 0.0276046, 0.1986246, -0.0285698, 0.0578464, -0.2685389, -0.0995264, 0.0299782, 0.3819751, -0.0731309, -0.0862887, 0.0655589, 0.1769768, 0.0374068, -0.0643319, -0.3037899, -0.2412053, -0.1300070, 0.0953529, 0.2455080, 0.1028997, 0.0496699, 0.2780990, 0.0436733, 0.0282080, 0.0183039, 0.0780210, 0.0553662, -0.0910214, 0.0227776, 0.1537467, -0.0238472, -0.1666262, -0.1455044, -0.0800281, 0.0998750, 0.4453037, -0.0928460, -0.0264877, -0.1433477, 0.0309958, -0.0464663, 0.0519355, 0.2386627, -0.0322981, 0.3918955, -0.1384275, -0.3730862, 0.1042562, -0.0840763, 0.1659195, -0.0741407, 0.0099414, 0.4528528, 0.0387757, 0.0270796, 0.1395009, -0.2743935, -0.1033302, 0.0350203, 0.1713298, 0.0308631, -0.0645609, 0.1552114, -0.0727325, 0.3354489, 0.0253301, 0.2735949, 0.1992740, 0.1817241, -0.1309627, 0.1303459, -0.0308000, 0.1408390, -0.0771936, 0.0268714, 0.0568418, 0.0408396, -0.0988570, 0.1019551, -0.0251061, 0.1617250, 0.3490078, -0.1046631, -0.0489336, -0.0358080, -0.1859378, 0.0085132, 0.1292803, -0.2492532, 0.1058178, -0.0184925, 0.0099441, 0.1682706, -0.0208473, 0.0147372, -0.0066501, -0.1781852, 0.0160379, 0.1589775, 0.0763847, 0.2812560, 0.2459783, 0.0687681, -0.0909406, 0.2519895, 0.2886911, -0.0103621, 0.1750779, 0.0305808, -0.3394182, 0.3790760, 0.2328954, 0.0304021, -0.1730505, 0.0849681, -0.0079131, 0.2168311, 0.0225064, 0.0612368, 0.0055914, -0.0283808, 0.3564338, -0.0637947, -0.1415868, -0.1191629, -0.0347170, -0.1001116, 0.2265013, 0.1521186, 0.2164169, -0.0102808, 0.3367968, 0.1525850, -0.0514733, -0.0946580, -0.0653857, -0.1149213, 0.0750685, -0.1537761, -0.1244465, -0.0909726, 0.1873952, -0.0913496, 0.0140599, 0.3778461, 0.1887102, 0.0570506, 0.2077320, 0.0450484, -0.1315451, 0.1800689, 0.1969139, 0.1246039, -0.0522698, 0.1531674, -0.2430759, 0.2572612, -0.1209005, 0.1529974, 0.0546396, -0.0258274, 0.4117777, -0.3743966, -0.0944431, -0.0516488, -0.0187969, 0.0104512, 0.1506363, 0.0501235, 0.1975297, 0.0969364, 0.2190267, 0.1809473, 0.0121413, -0.0469255, -0.0677327, -0.0919020, 0.0523575, -0.1166499, 0.0131582, 0.0016223, 0.1828314, 0.0317480, -0.0603651, 0.0168355, 0.2381065, -0.0644196, 0.1214829, -0.1402263, -0.2580840, 0.2939126, 0.0929884, -0.1482369, -0.0562798, -0.0159296, 0.0063701, 0.1752317, -0.1051414, 0.0065816, 0.0306327, -0.0749477, 0.1573239, 0.0090140, 0.0458717, -0.2257026, 0.0134158, -0.0121276, 0.3021936, 0.1447391, 0.0198012, 0.1730571, 0.2748802, 0.0280657, -0.0085231, -0.2373109, -0.0838828, -0.0626611, 0.0546418, -0.0273715, 0.0127199, -0.1693058, 0.1465559, -0.1347251, 0.1167072, 0.0554091, 0.1067030, 0.0289027, -0.0101264, -0.0062137, 0.0952583, 0.0900537, -0.0854528, -0.0488368, -0.0036252, 0.1682309, 0.4211317, -0.1011828, 0.0762080, -0.0247690, 0.0836274, 0.0448115, -0.1566464, 0.2131029, 0.1210317, 0.2324871, -0.1040523, -0.2412765, 0.0562330, 0.0053879, 0.0016889, 0.0103561, 0.0836141, 0.2372961, 0.0746417, 0.1163326, 0.0532555, -0.1486807, 0.0255499, 0.0501690, 0.0058099, -0.0037226, -0.0151310, 0.0382395, -0.1771977, -0.1179370, 0.0291547, 0.0565185, 0.2065892, -0.1283626, -0.0317070, 0.1043827, -0.0804745, -0.0451716, 0.0454750, 0.0303341, -0.1094946, 0.0717386, -0.1339175, -0.0882287, 0.0072388, -0.0070601, 0.1199960, -0.0395891, 0.0799698, -0.1183696, 0.1843316, 0.0461558, 0.1383476, 0.1011766, -0.1026275, 0.0384017, 0.0244378, -0.1866957, 0.0694735, -0.0862908, -0.0977887, 0.0720473, 0.0843523, 0.0535606, 0.1790757, 0.0385843, 0.1664081, -0.0886817, 0.0540752, 0.2024199, 0.2969318, 0.1360566, 0.2640443, 0.0612300, -0.3711911, 0.5722917, 0.1883611, -0.1091309, 0.0160806, -0.1278029, -0.0727495, 0.3697583, -0.0863324, -0.0354410, -0.0324638, -0.0513397, 0.3496298, -0.0780670, 0.0964050, -0.2918820, 0.0476868, 0.0051698, 0.4891298, 0.2158738, 0.0497583, 0.3254720, 0.3068710, 0.0568265, 0.0998509, -0.2681111, -0.2179232, -0.0594104, 0.0861655, 0.1221441, 0.0927776, -0.1812803, 0.3288058, -0.1350615, 0.1249707, -0.0480614, 0.0099242, 0.0108524, 0.2002075, -0.0155853, -0.0771127, 0.0106385, -0.1144631, 0.0938256, 0.1099462, 0.0262388, -0.0417353, 0.0406899, 0.1173594, 0.0557942, 0.0209506, 0.1241499, 0.0149975, -0.0231014, 0.0549717, -0.1268896, 0.2155925, 0.1586458, 0.0339958, 0.1837280, -0.1115026, 0.1317426, 0.0544162, -0.1891286, 0.0968895, -0.0773559, -0.0006247, 0.2329849, 0.2522520, 0.1340773, -0.0262505, -0.0110373, 0.1586221, -0.2438082, 0.0907695, -0.0068979, -0.0756581, 0.1525604, 0.1498764, 0.0792192, 0.0727572, -0.0950013, 0.0458045, 0.0532070, 0.0376727, -0.1181954, -0.0515692, -0.0514270, -0.0642803, 0.0075158, -0.2537528, 0.0550820, 0.0086680, 0.1020255, -0.0384035, -0.0296152, -0.0739848, 0.1157653, 0.1282831, -0.1494079, -0.3352095, -0.1855527, -0.1174976, -0.1021687, -0.1195255, -0.2581396, 0.1161277, 0.0687329, 0.1218027, 0.3023509, -0.0423620, 0.2672545, 0.2212545, 0.0567080, 0.1280476, 0.0034356, 0.1692715, -0.0186707, -0.2514981, -0.0421485, 0.1070573, 0.0454740, 0.0814534, -0.0253220, -0.1064432, 0.0386227, 0.4243780, 0.0673514, 0.0445206, -0.2274008, -0.0689689, -0.1269779, 0.0947194, 0.2739683, -0.0414276, 0.2207769, -0.1652095, -0.3207724, 0.0756820, -0.1800167, 0.1341016, -0.1277603, 0.1118644, 0.2531807, -0.0239171, 0.0416604, 0.1836447, -0.2280639, -0.4259863, 0.0431790, 0.2325373, 0.0522770, -0.3137045, 0.1898074, -0.0283242, 0.5136158, -0.0526263, 0.3134669, 0.0827940, 0.4331023, -0.2785960, 0.2378170, -0.1718848, 0.2840393, -0.0738651, 0.1276468, 0.0491142, 0.0724916, 0.0944150, 0.1615584, 0.0187391, 0.5009721, 0.3165060, -0.3028131, -0.0450312, 0.0030985, 0.2708218, 0.1690821, -0.1586524, -0.1752167, 0.1579420, 0.1023560, -0.0245807, 0.1536802, -0.1976039, -0.1003954, 0.0508191, -0.0079922, -0.0075539, -0.0425409, 0.1197831, 0.1056905, 0.0844729, -0.2120419, -0.2671377, -0.4136035, 0.2558374, -0.0805482, 0.0975428, -0.4411223, 0.0866302, 0.2218378, 0.1889997, 0.0344980, 0.0631849, -0.0908859, 0.0463600, 0.1447899, 0.0934084, -0.0793260, -0.2206043, -0.1738649, -0.0030359, 0.3036871, -0.0569196, -0.1382490, -0.0315118, 0.1163319, 0.1098552, 0.1931170, -0.1331010, -0.0662209, 0.1373620, -0.0416974, -0.1841499, -0.2297016, 0.4867609, 0.1408280, -0.1419996, 0.1164926, -0.1169445, 0.1792517, 0.0997180, -0.0930852, 0.2665899, 0.1772826, 0.2911820, 0.0544398, -0.0070780, 0.0365776, 0.0129455, 0.0703210, 0.1501381, -0.0386450, 0.0326638, 0.1565036, -0.1359735, 0.1759621, -0.0549826, 0.1268574, 0.1616875, 0.0543186, 0.0347628, -0.1171480, 0.1026899, 0.0547493, -0.0986320, -0.1110825, -0.0390160, 0.0535269, 0.1375834, -0.0075321, 0.2022396, 0.3148380, 0.0665971, 0.1468842, -0.0530879, -0.0454508, 0.0529535, -0.1947910, 0.0460920, -0.1431887, 0.0155312, 0.1224896, -0.0673204, -0.2217153, 0.0917101, -0.0985135, 0.0458894, -0.1854495, 0.0945850, 0.1473071, 0.1370154, 0.0041797, 0.1359116, -0.0341140, -0.0019052, 0.1315651, 0.0324863, 0.0002158, -0.0819791, -0.1324055, 0.0687811, 0.1051465, -0.0008062, -0.1634116, 0.0080519, 0.0435474, 0.1111137, 0.1583468, -0.3895085, 0.0376045, 0.0552615, -0.0420488, -0.0292832, -0.1793548, 0.1940987, 0.0951184, -0.0234378, 0.0835786, -0.0221211, 0.0981485, 0.0474826, -0.0427655, 0.2057450, -0.0600090, -0.1011127, -0.0368723, 0.1319060, 0.0708340, 0.2680511, -0.0411812, -0.3372578, -0.0255649, 0.0765969, 0.1671286, 0.2167058, -0.1751426, 0.2182699, 0.0899920, -0.0033912, 0.0165648, -0.2012881, 0.3050904, 0.0641010, 0.2143210, 0.0976318, 0.0817550, 0.1798538, 0.2406318, -0.1867285, 0.0467752, -0.2025434, 0.0962502, 0.2255851, 0.0721069, 0.0202640, 0.0537253, 0.2397274, 0.2431281, -0.1201723, 0.1241195, 0.1453437, -0.1557724, -0.1263190, 0.2886108, -0.0805936, 0.2567955, 0.1924004, 0.1736066, -0.1675311, 0.1188851, -0.1315535, 0.1202336, -0.1623448, 0.0034862, 0.0011807, -0.0605923, -0.1432793, -0.0043426, -0.1146239, 0.2328805, 0.3920560, -0.1398847, -0.0989397, -0.1441049, 0.1094199, 0.1353636, -0.0342076, -0.1263096, 0.0920982, -0.0223685, 0.0073325, 0.1180372, -0.2517564, -0.3154455, 0.0648174, -0.0863338, -0.0438278, -0.0120813, 0.1211038, 0.1419234, 0.2247398, -0.1210846, 0.0668434, 0.0613511, -0.0599937, 0.1244880, 0.0679014, 0.0169780, 0.0859863, -0.0299121, 0.0579265, 0.1274457, 0.1369797, -0.0142882, -0.0152089, 0.1057995, 0.0139639, 0.0978561, -0.1101636, 0.0624334, 0.3387574, 0.0274576, -0.0464072, 0.0565576, 0.0334890, 0.2432028, 0.1288034, -0.0277457, -0.0693631, -0.0557014, -0.0787942, 0.0252883, -0.0541283, -0.0581677, 0.1166344, 0.1466553, 0.0611536, 0.1517839, 0.1539167, 0.1629883, 0.1395402, 0.1281774, 0.2036290, 0.0583166, 0.1824410, 0.3300922, 0.2729586, 0.0368477, -0.0773251, 0.1297181, -0.2295886, 0.1342872, -0.1510844, 0.1567210, 0.0914983, 0.0273497, -0.0945633, 0.0131086, -0.0095299, 0.2521878, 0.2160577, -0.0042421, -0.0637379, -0.1271943, 0.1970858, 0.1724376, -0.0199014, -0.0019749, -0.0008311, 0.0532547, 0.1517689, 0.0165826, -0.0869183, -0.2509376, 0.1268211, 0.0040535, 0.1554221, 0.0672799, 0.0776693, 0.1677678, 0.3528205, -0.3164931, 0.0200708, -0.1696217, -0.0048509, -0.0180708, 0.0915937, -0.0282529, 0.0483110, 0.1751201, 0.0456137, -0.2793117, 0.0869260, 0.0756640, -0.0060428, -0.0244918, 0.0556037, -0.0454325, 0.0620784, 0.0531370, 0.0376116, -0.0324388, 0.2129904, 0.0474446, 0.2094311, 0.0709239, 0.0563645, 0.0939073, -0.0209472, 0.2123675, -0.0040568, -0.0202855, 0.1694612, 0.0818217, -0.0133929, 0.1541006, 0.0609884, -0.0297489, 0.0877483, -0.1948574, 0.1109802, -0.0141827, 0.0719839, 0.1544085, 0.0651931, -0.1164017, -0.3476659, 0.0671368, -0.0120933, 0.3118630, 0.4476832, 0.2477911, -0.0374006, 0.1289403, 0.3391702, 0.1810415, 0.4087949, 0.0255976, -0.3636750, -0.0277944, 0.2770663, -0.0858706, -0.2039078, 0.0640655, 0.1046631, -0.0790921, -0.1587275, -0.3282816, 0.3149728, 0.2542259, 0.1789556, 0.2293674, -0.1377006, -0.1724912, 0.4153343, -0.0533522, -0.3121149, -0.0342609, -0.0364869, 0.3173378, -0.2527095, 0.0227176, 0.1241251, 0.4643567, -0.2299815, 0.1643298, -0.0419958, 0.5448251, -0.2439101, 0.2388859, -0.3929267, 0.2709555, 0.0788806, -0.0731085, 0.1819758, -0.1043447, 0.2842651, 0.1419394, -0.0517220, 0.2201522, 0.2309805, -0.2302336, -0.0345637, 0.0133205, 0.2205119, 0.1287036, -0.1604019, -0.1039510, 0.0815864, 0.1784894, -0.1448413, 0.0313534, -0.0937422, 0.0175420, 0.0904810, -0.0706644, 0.0103337, 0.1057760, 0.1232812, 0.2231040, -0.0929260, -0.0224973, -0.2216284, -0.2759682, 0.1242518, -0.2273744, -0.0851852, -0.4107179, 0.2830814, -0.0573786, 0.2900250, 0.0703388, 0.2367309, -0.0353033, -0.0461389, 0.0757540, -0.2633409, 0.0834944, -0.1310984, -0.3587838, 0.3628905, 0.0782126, -0.2231306, -0.1888587, -0.0545586, 0.2527952, -0.1067689, -0.0064214, 0.2578904, -0.2258448, 0.0445774, -0.0373641, -0.1511404, -0.3211170, 0.5739539, 0.2382930, -0.2092171, -0.1156397, 0.0843561, 0.3120153, -0.0954690, 0.1854065, 0.3495750, -0.1736812, 0.2365922, 0.0692179, -0.0990338, -0.1231851, 0.2150815, -0.1306803, 0.1156135, 0.0162113, 0.0349834, 0.0406373, 0.2131620, -0.0459964, -0.0649705, -0.0143496, -0.0190454, 0.0097475, -0.0655613, 0.2747841, 0.0043188, 0.1191312, -0.0779188, -0.0143105, -0.1296676, -0.0674693, -0.1245580, -0.1032700, 0.0586838, -0.0287370, -0.0903502, 0.0179240, 0.2929253, 0.0547910, -0.1412193, -0.0148449, 0.0636778, 0.0896431, -0.0885704, 0.0818911, 0.1182231, -0.4259281, 0.1019717, -0.3549793, 0.0385020, -0.5459166, 0.2702778, 0.0308811, 0.1369698, -0.0535592, 0.1112488, 0.0676692, -0.0578505, 0.1180220, -0.1704092, 0.0052057, -0.0725868, -0.2203720, 0.1938023, 0.1353357, -0.1081495, -0.1874768, -0.0424991, 0.1919333, 0.1097804, 0.1999698, -0.0964925, -0.1249383, 0.0099438, 0.0204972, 0.0186865, -0.2196877, 0.2100696, 0.2370404, -0.0340972, -0.0862417, -0.0841479, 0.1292686, 0.0762949, 0.0959898, 0.3140408, -0.4084839, 0.0740187, -0.4006624, 0.0846595, -0.2030533, 0.3111199, -0.0645724, -0.3006584, -0.0081231, 0.2087855, 0.1776381, 0.1702383, 0.0036760, 0.2831955, -0.0147580, -0.0652945, -0.1196921, -0.2686384, 0.3258738, 0.0405119, 0.1082629, 0.1155132, 0.1221959, 0.2071721, 0.7456440, -0.2682689, 0.0498060, -0.0539512, -0.0458301, 0.0914590, -0.0568602, 0.1222316, 0.2177871, 0.2081797, 0.2643073, -0.3640482, 0.1304058, 0.0794319, -0.2636914, 0.0714720, 0.3038584, -0.0878149, 0.1689495, 0.0831233, 0.3947182, -0.2278300, 0.1854807, -0.5335009, 0.0885407, -0.0189534, -0.1619901, 0.1775887, -0.3098898, 0.0680178, 0.0066493, -0.1724831, 0.1547397, 0.1921853, -0.0100354, -0.0225388, -0.0482945, 0.0034749, 0.0873296, 0.0768844, -0.2345435, 0.0696113, 0.0842791, 0.0012031, -0.0759819, -0.1424875, -0.0509689, -0.0752677, -0.2686817, 0.0280172, 0.2515833, 0.0468994, 0.0954919, 0.0472130, 0.0118068, -0.0840062, 0.3757174, -0.1149149, -0.0351747, -0.1133074, 0.3945434, -0.0945029, 0.0891566, -0.1022894, 0.1489211, 0.3598934, 0.0228314, -0.0902228, -0.0283526, 0.2842809, 0.3012520, 0.1423986, 0.1530422, 0.0763298, -0.2662569, 0.5281415, 0.2439428, 0.1649843, 0.2768130, 0.0223604, 0.0868692, 0.1026028, 0.3543645, 0.0105140, -0.1248850, 0.3400951, 0.3535477, -0.2195097, 0.1874961, 0.2248434, 0.0500370, 0.0958707, -0.2496917, -0.1939913, 0.1366424, -0.0815197, 0.1819752, 0.0824174, 0.1507705, 0.1191345, 0.2654988, -0.2312119, 0.1361166, -0.1956506, 0.1250602, -0.0278156, -0.1684859, 0.0956496, -0.1466562, 0.0653168, 0.0644698, -0.0924969, 0.1579335, 0.1545208, -0.0205970, 0.0648629, -0.0373382, 0.0368595, 0.1531642, 0.1060842, -0.2268278, -0.0112675, 0.0930384, 0.1789942, -0.0906527, -0.0819785, -0.0107448, -0.0789668, -0.1863945, 0.1057726, 0.2891479, 0.1155242, 0.0114967, 0.1069884, -0.0117348, -0.0069406, -0.2553782, 0.0038099, 0.0552232, 0.0175569, 0.0028230, 0.1068024, -0.1100429, -0.0318050, -0.0415117, 0.0697467, -0.0254069, -0.0468472, -0.0777797, -0.0240773, 0.0084114, 0.0405372, 0.0358030, -0.0849677, 0.0903276, 0.1726640, 0.0116666, 0.0544490, 0.0877725, -0.0391104, 0.0125117, -0.3949948, -0.0079627, 0.0226369, -0.2536785, -0.0249237, 0.0585688, 0.0140999, 0.1253929, 0.0119074, 0.0551289, 0.0762838, -0.0477681, 0.0324982, 0.0288493, 0.0919705, 0.3779339, -0.3331796, 0.2007893, -0.1726793, 0.5365922, -0.0585332, 0.0917568, -0.2471654, 0.4183583, -0.0250867, 0.4007334, 0.3202589, -0.1855118, 0.5002189, 0.0818017, 0.0673225, 0.2819993, 0.2582466, -0.0986213, -0.0974056, 0.4149181, 0.4479879, 0.2100879, -0.2593095, -0.0393042, 0.2098121, 0.2821132, -0.2381986, 0.2351533, 0.0217529, 0.0736737, 0.3033642, 0.0505228, 0.0491839, -0.1403535, 0.0412747, 0.1855997, -0.2884952, -0.0575630, -0.2199185, 0.3169606, -0.0743003, 0.1060511, -0.1460739, 0.2673158, -0.1374191, 0.1182191, -0.2918414, 0.1811889, -0.1114185, 0.0945262, 0.1792995, -0.1372634, 0.2621058, 0.0318214, -0.0391163, 0.2022329, 0.0026963, -0.0110412, -0.1304135, 0.1402300, 0.1479346, -0.0286170, -0.1385071, -0.0617535, 0.0846403, 0.1224038, 0.0004866, 0.1808242, -0.0396092, 0.0283209, -0.0523378, -0.1815699, -0.0081625, -0.0673563, 0.0064328, 0.1610001, -0.0960691, -0.1997841, -0.3198293, 0.1522148, -0.0257744, -0.0226474, 0.1623929, 0.0631538, -0.1503823, 0.3214246, 0.1211633, 0.1859556, 0.1707723, 0.1144571, -0.0377355, 0.1814972, 0.1671701, 0.1989699, 0.1032160, 0.0020528, 0.1553799, -0.3062166, 0.1197483, -0.1153034, 0.3516244, 0.1026282, 0.0906545, 0.3324026, 0.0698252, 0.3918035, 0.1211530, -0.0036834, 0.0342929, -0.0726243, 0.1347301, 0.1050123, 0.1918691, -0.1413158, 0.1031597, -0.0688241, -0.0122070, -0.2015107, 0.0733609, -0.1282799, -0.0210960, -0.0895506, -0.0170459, -0.1910985, 0.3763955, -0.2723860, 0.3008282, 0.2168916, 0.2398573, 0.0853637, -0.1198472, 0.0267400, -0.1208313, 0.3994486, 0.0128937, -0.1606963, 0.1884048, 0.0167639, -0.1357943, -0.1036241, -0.2360173, 0.2838593, -0.1723818, -0.0134910, 0.1047089, -0.2556389, 0.0431921, -0.1318795, -0.1565483, -0.1458418, 0.3049258, 0.2150912, -0.1208631, -0.1072938, -0.1349450, 0.3395818, -0.0172538, 0.2680461, 0.2662638, -0.4970317, 0.1538017, -0.2266079, 0.4554995, -0.4030932, 0.0241911, 0.3630141, -0.1508763, -0.3052724, 0.1305191, 0.1537001, 0.1171078, 0.0244289, -0.0834728, -0.4534850, -0.1481970, -0.2346289, 0.0978074, 0.1603136, 0.2281485, -0.1086829, 0.3007004, -0.0460775, 0.5789331, 0.6387429, -0.2287703, 0.3714036, 0.0218829, 0.1593084, 0.1754071, -0.2266179, 0.2793485, 0.1976435, 0.2893304, 0.4635845, 0.2819348, -0.0835880, 0.4406214, -0.1838998, 0.2153038, -0.3992608, 0.0408452, -0.3936059, 0.1305479, -0.3631929, 0.1134881, -0.0211070, -0.1440576, -0.2374878, 0.1090502, 0.0392677, 0.0083447, 0.1212540, 0.0313217, -0.1072166, 0.0513591, -0.1534570, -0.1544561, 0.2039653, 0.0855184, -0.0951758, 0.0643879, 0.0968248, 0.4299633, 0.5424745, -0.3717279, 0.0553645, 0.0099891, 0.0332046, 0.1879375, -0.1545957, 0.1316505, 0.2058910, 0.1671457, 0.1803628, -0.0127131, 0.0300194, 0.0984607, -0.1269942, 0.1735023, 0.1688373, 0.0808166, 0.0298312, 0.0869670, 0.1261673, -0.1729414, 0.0878988, -0.3493914, -0.0695719, -0.0874117, -0.0554185, 0.1277231, 0.1021345, 0.2111150, -0.1764307, -0.1417039, 0.0180583, -0.0457616, 0.1277621, -0.0703545, 0.1015398, 0.0496272, -0.1550216, 0.2590737, 0.0159401, 0.0361908, 0.1594941, 0.0149759, 0.0358684, 0.0096461, -0.0450648, -0.0840731, -0.1866910, 0.0920185, 0.3141201, -0.0784492, 0.0602430, 0.1381536, -0.1915216, -0.1360847, 0.2910327, 0.0166257, -0.1772997, -0.0425941, 0.3005095, -0.0775231, -0.0266582, -0.0230048, 0.0872576, 0.1819755, -0.0018982, 0.0276334, 0.0565216, 0.2828892, 0.2199281, 0.1254633, 0.0268731, -0.1050830, -0.0093827, 0.1723511, 0.3085960, 0.1135140, -0.0175422, 0.0254729, 0.1801013, 0.0814893, 0.2312442, -0.0419373, -0.0670168, 0.2536175, 0.1619502, -0.2468528, 0.0604604, 0.2776412, 0.0057474, -0.0908495, -0.0875275, -0.1451850, -0.0228111, -0.1765662, 0.1057382, 0.1241332, 0.0128148, 0.1217481, 0.1804959, -0.1309088, -0.0308060, -0.0415266, 0.1021474, 0.0147159, -0.0659484, 0.0154524, 0.0509109, 0.1473719, 0.1367746, 0.0049268, 0.0989094, 0.0772387, 0.1431008, 0.0192590, 0.0381420, -0.0989385, 0.0673607, 0.0374940, -0.0169531, 0.0179956, 0.0339629, 0.0318401, -0.0450840, 0.0108838, 0.0186030, -0.0814650, -0.0536074, 0.1195013, 0.2224859, -0.1554033, 0.1043000, 0.1490091, -0.0396010, -0.0207322, -0.0668252, -0.0285929, -0.0461695, -0.0439064, -0.0359442, 0.0533210, -0.3033175, 0.0626940, 0.0903523, 0.0599859, 0.0165022, -0.0672648, -0.0482395, -0.0252578, 0.2097165, 0.1734049, 0.0748091, 0.0606162, 0.0069681, -0.0762280, -0.0267916, -0.0255343, 0.2647512, -0.0617531, 0.0099262, -0.2446314, -0.1495145, 0.0735983, -0.1848365, -0.0489289, -0.0131526, -0.0322198, 0.1344172, 0.0704069, -0.0376958, -0.1835543, 0.1590182, 0.0014058, -0.0159551, 0.0563825, 0.1496891, -0.0542694, 0.1162410, -0.0467994, 0.2380764, 0.1795036, -0.0374526, -0.3408541, 0.1773441, -0.0778227, 0.6624670, 0.2856180, -0.2222566, 0.3890345, 0.0779408, 0.1515224, 0.2860934, -0.1532074, 0.1368199, -0.0075336, 0.4929797, 0.4693128, 0.0642076, -0.1484178, 0.2134319, 0.1153041, 0.2277015, -0.1204014, 0.3150825, 0.1983345, 0.0550845, 0.1230248, 0.2284103, 0.2597835, -0.2540803, 0.1201588, 0.0781178, -0.1477641, -0.0991390, -0.2466474, 0.1123410, -0.1256617, -0.0155707, 0.0891706, 0.0976188, -0.0387359, 0.1823566, -0.1092074, -0.0090315, 0.0702712, 0.0594849, 0.0792025, -0.0342215, 0.1746882, -0.1518261, -0.0938948, -0.0271978, 0.0938307, -0.0963615, 0.0077476, 0.1205111, 0.1870723, -0.0423720, 0.0465713, 0.0800419, 0.0821748, 0.2263056, -0.1131474, 0.1532576, 0.1106299, -0.0106807, 0.0242833, 0.0637727, 0.0645515, 0.0554729, 0.1373807, 0.1014390, 0.0484578, -0.0835293, -0.0283346, 0.1585160, 0.0286567, -0.2804472, -0.0606013, 0.1467351, -0.1410394, 0.0611486, 0.1535671, -0.0800921, 0.2714658, -0.0601713, -0.0570389, 0.0211810, 0.0839924, 0.0907233, 0.0856400, 0.0038868, 0.2353165, 0.0043589, 0.2820182, 0.0699790, 0.0261533, 0.0576866, 0.1559366, 0.2162789, 0.0118956, 0.2227638, 0.0606465, -0.0663127, 0.2711236, 0.2290319, -0.1846901, 0.1659428, 0.0773437, -0.0454417, -0.1064762, -0.2224667, 0.0065115, -0.0051188, 0.1076582, 0.3014049, -0.0313995, 0.1589174, 0.3138995, 0.2649204, -0.0130472, 0.3195731, -0.0390334, 0.0126609, 0.0898037, -0.0899293, 0.1347037, 0.0131423, 0.0564530, -0.1241802, -0.0787482, 0.0625769, 0.4225606, 0.2279718, 0.1078063, 0.1945599, -0.0018825, -0.0414232, 0.3670290, 0.0707412, 0.2672088, 0.2481320, 0.0126231, 0.2636248, 0.2179081, 0.0407740, 0.0221425, -0.1614270, 0.1173745, 0.3290016, 0.1664982, 0.0858370, 0.2123957, 0.0817211, -0.0212251, -0.0005551, 0.1493842, -0.1624763, 0.0282145, 0.0214730, -0.0569945, 0.0869176, 0.1993899, -0.0862246, 0.1040314, 0.0431894, 0.2668693, 0.0954544, 0.4356057, -0.0635643, -0.0790145, -0.0981650, -0.1188299, 0.3077695, 0.0142526, 0.1172816, -0.0320687, -0.0028560, 0.1721650, 0.3366380, 0.0054901, 0.0124590, 0.1595554, 0.0166998, 0.1732469, 0.0176942, 0.1980539, -0.0816261, 0.1206813, 0.2280039, -0.1878292, -0.0117586, 0.0424355, -0.0562982, 0.0539031, 0.0016639, 0.0175611, 0.0539848, 0.2335620, -0.0163350, 0.2241043, -0.0211916, -0.1026794, 0.0349034, -0.1652614, 0.1864364, 0.2034337, -0.0659805, 0.1438320, -0.3160794, -0.2048448, -0.0180279, -0.0447578, 0.1666442, -0.0342967, 0.0766209, 0.0525764, -0.0857177, 0.2826692, 0.2107199, 0.0389231, -0.0797000, -0.0093641, 0.2184675, 0.1723681, -0.0230925, 0.2416588, -0.0209176, 0.1826027, 0.2022525, 0.0177556, 0.2987073, 0.2481931, -0.1102722, -0.1167044, 0.0160351, -0.0820093, -0.0615353, 0.1278675, -0.0273395, -0.2543565, 0.2960419, -0.1472568, -0.0295665, -0.0898276, 0.0055736, 0.0829042, 0.0473162, 0.0752161, -0.3565159, -0.1265212, -0.0111110, -0.0306755, -0.0445523, -0.0216494, -0.0531430, 0.1727236, -0.1038673, 0.2440962, 0.2747497, 0.0484549, 0.3496753, 0.0056224, 0.0694921, 0.0804773, -0.1132254, -0.0216479, 0.0005220, -0.0040859, 0.1536831, 0.0495742, -0.1221322, 0.0663005, -0.2256109, -0.1397598, -0.0751490, -0.0957104, 0.0072429, 0.0825280, -0.0539534, 0.1566175, -0.1313618, 0.0596027, 0.0307440, 0.0925107, -0.1264466, -0.1359149, -0.2049449, -0.1911218, 0.0519601, -0.0326971, -0.0716721, 0.0329923, 0.0701965, -0.0010436, -0.0612618, 0.0462665, 0.1182863, 0.0132833, -0.0536650, -0.0756561, -0.0157820, -0.1341165, -0.1584192, 0.0600668, -0.0739695, 0.1277794, 0.0727160, 0.0501449, 0.0477353, 0.0699452, 0.0934274, 0.0769574, 0.1150260, 0.0599445, 0.0943615, -0.2111203, -0.0444885, -0.0601772, 0.0830781, -0.0913955, 0.1379317, -0.0946652, -0.0316969, 0.1088738, 0.0818273, -0.0789403, -0.1121935, 0.1419611, -0.0932568, 0.0222821, 0.0115548, -0.0591928, -0.1688217, 0.0507436, 0.1165169, 0.2657143, -0.0143101, 0.0162930, 0.0582716, -0.0594479, 0.3476352, -0.1475322, -0.0715088, 0.1446379, 0.0484287, -0.0318070, 0.0657187, 0.0136161, 0.0278033, 0.1545877, -0.0592786, -0.0378826, -0.0741290, -0.1797023, -0.0584931, -0.0868086, -0.1632000, 0.0977491, 0.0297982, 0.2325948, -0.0137758, 0.1165432, 0.0737304, 0.3581679, 0.1040542, -0.2461189, -0.0952825, -0.0732346, 0.1889021, 0.2365600, 0.0725396, 0.0801036, -0.2433263, 0.1973117, 0.0845352, 0.2828246, 0.2213288, 0.0842379, 0.2239240, -0.2209137, 0.2538530, -0.1502572, -0.1711968, 0.2559465, 0.0886124, -0.0592338, 0.3019627, 0.1746448, 0.0543442, 0.1529985, -0.0986306, 0.1644742, -0.0345814, 0.1523341, -0.0114726, 0.0644708, 0.0600256, 0.0791032, -0.0312498, 0.0736796, -0.0430327, -0.0562159, 0.0251398, -0.1136785, 0.0220870, -0.0420634, -0.1022629, -0.0381456, -0.1016117, -0.0337885, -0.0086374, -0.0331742, 0.1243683, -0.1634357, 0.0066130, -0.0605105, -0.1633413, -0.0173947, -0.0284350, 0.0730683, -0.1518236, -0.0098218, 0.0885277, 0.0748884, -0.0936240, 0.1729562, -0.0967456, 0.0027524, 0.0327044, 0.0653295, 0.0717818, 0.0705097, -0.0077875, 0.0092109, 0.0489954, 0.0283550, -0.0424663, -0.0587633, 0.0302622, -0.1551957, 0.2883229, -0.3735371, -0.0319596, 0.1235673, 0.0319965, 0.1142806, 0.0853927, 0.2021170, -0.1654835, 0.0347479, 0.0253620, 0.0717602, -0.0498954, 0.2408537, -0.0072512, 0.1920467, -0.0353376, 0.1403110, 0.1748656, 0.0834756, 0.4724808, 0.1389830, -0.0366417, -0.0197263, -0.0036474, 0.0041942, 0.0628797, -0.0981734, 0.1173345, 0.1220539, -0.0634993, -0.1134647, -0.0755313, 0.0400450, -0.0151675, 0.2287636, -0.1943709, -0.1317284, -0.0328366, -0.0768794, 0.1929236, 0.2403952, 0.0845221, 0.4107741, -0.2704249, 0.0320627, 0.2056496, 0.1795227, 0.2914478, -0.1524897, -0.2262623, 0.3213210, 0.1358803, 0.0613863, -0.2432298, -0.3602407, 0.1060914, 0.0360312, -0.0399945, 0.3255664, -0.0046390, 0.3174735, -0.1251500, -0.0106545, -0.0988853, 0.2488076, 0.1037145, -0.1100697, 0.2740440, -0.2242421, 0.1190877, -0.0614087, 0.1180410, 0.3177331, 0.2251695, -0.0967520, -0.0736613, -0.0880474, 0.2135104, 0.1619440, 0.1121995, 0.0991702, 0.0499477, 0.1499362, -0.2582387, 0.2422641, -0.1007862, 0.1248454, 0.0798230, -0.3493113, -0.1843482, 0.6873617, -0.0015148, -0.1559610, 0.2586505, -0.4841425, 0.0026527, 0.3362826, -0.4844767, 0.6771153, -0.0182661, -0.0451828, 0.3245613, 0.0783477, 0.2050133, 0.1888837, -0.1794487, -0.2421736, 0.2202877, -0.0538566, 0.3917046, 0.0462903, 0.5143296, 0.0008751, -0.0135002, 0.0624296, -0.1535297, 0.0852108, -0.0141296, -0.1052564, 0.1316494, 0.0979113, 0.0626237, 0.0543732, 0.0437085, 0.3084924, 0.1054642, 0.2715148, -0.1109071, -0.1586413, -0.1223051, -0.0161536, 0.0628282, -0.1055928, 0.0822015, 0.0573507, -0.1080897, 0.0597405, 0.0792483, 0.0259985, 0.0594393, -0.0222393, 0.1640731, 0.1326687, -0.0792401, 0.1743508, -0.0326227, 0.0127271, 0.0517678, -0.0930289, 0.0452359, 0.0619075, -0.1511738, 0.0317377, -0.0643779, 0.1687538, 0.1527865, -0.0158982, -0.0520989, 0.1570354, 0.0060550, -0.3031828, -0.1812776, -0.1211455, 0.1078257, 0.1469245, -0.0336818, -0.0620995, -0.3181101, 0.1717681, 0.0654248, -0.1259069, 0.1058671, 0.0896540, 0.0551866, -0.0972993, -0.1893384, 0.0632741, -0.0108594, -0.0194192, -0.0371084, 0.1613375, 0.1007414, -0.0367399, 0.0665431, 0.1202008, -0.1026210, -0.0560626, -0.0354040, 0.0888368, -0.0013581, 0.0229435, 0.1341169, 0.0877135, 0.0806891, 0.0642451, -0.0716569, 0.1226181, 0.0037502, -0.2698954, 0.2270379, -0.0987777, -0.0632531, 0.0023417, -0.0953645, 0.1145498, 0.1294708, 0.0598387, -0.2379022, -0.1385108, -0.1277252, 0.0195173, 0.0143290, 0.0276562, -0.1278231, 0.0929973, -0.0434191, 0.1291679, 0.1399277, 0.0234037, 0.2540445, 0.0119292, 0.0637979, 0.0109945, -0.1004908, -0.0223922, -0.0244899, -0.0177171, 0.0143478, 0.0101488, -0.0705593, 0.0543904, -0.1221263, -0.0238939, -0.1075226, -0.0797634, 0.1080424, 0.2467884, -0.0603431, 0.1399801, -0.2457328, 0.1124367, 0.1424566, 0.1788162, -0.0976078, -0.2887048, -0.0837905, -0.2914831, 0.1154264, 0.0074982, 0.1090475, -0.0482388, -0.1119784, 0.1195390, -0.0766293, 0.1628080, 0.2514575, 0.0225955, 0.0155967, -0.4772575, -0.0561108, -0.1191893, -0.2404904, 0.0298594, -0.0255122, -0.0039506, 0.2870604, 0.2886504, 0.1130757, 0.0253133, 0.0981089, 0.3224015, 0.0717274, 0.2192709, 0.1353867, -0.1065955, 0.0126273, -0.1045549, 0.1496995, -0.0914439, 0.1507616, -0.2736477, 0.0451098, 0.0557284, 0.2331562, -0.1078961, -0.0844879, 0.2552190, 0.0476150, 0.1556284, 0.1556779, 0.1086294, -0.1506194, 0.1376749, 0.2116242, 0.2375878, 0.0623757, -0.0416863, 0.1544701, 0.0644935, 0.3458113, -0.0772180, -0.0937625, 0.0882296, 0.0917221, 0.0425767, 0.1957248, 0.0756053, -0.0899542, 0.1185128, -0.1414025, -0.1213748, -0.0692685, -0.0633835, -0.0977665, 0.1143807, -0.3759568, 0.2653197, -0.0195834, -0.1195500, -0.0195894, 0.1131777, 0.0856336, 0.5092497, 0.1636985, -0.3319544, 0.0697216, -0.0994075, 0.2248232, 0.2141164, 0.1842617, -0.0619714, -0.1414582, 0.4741428, -0.0070904, 0.4321566, 0.3125622, 0.0771746, 0.5019433, -0.3854191, 0.3456171, 0.1056829, -0.3369399, 0.2998368, 0.0739064, -0.3017284, 0.4573635, 0.4184372, 0.0937922, 0.0141937, -0.3288351, 0.1844924, -0.2209341, 0.2386007, -0.0726642, 0.1073994, 0.0386609, 0.0008513, 0.0185482, 0.0383128, -0.0570663, -0.2283143, -0.0680107, -0.1009854, 0.0029615, 0.0707595, -0.2076246, -0.0204342, -0.2096528, -0.0494032, 0.0198837, -0.1504729, 0.0925548, -0.0327424, 0.0060573, -0.0740985, -0.1465689, 0.0361967, -0.0922875, -0.0780784, -0.0973841, 0.0014753, 0.0091809, 0.0048044, 0.0277445, 0.0717318, -0.1122698, -0.0488855, 0.0328702, 0.0360227, 0.0179612, 0.0640182, 0.0588300, -0.0134582, 0.0423927, 0.1936332, -0.0405882, -0.0432564, 0.0088989, -0.2396587, 0.3350563, -0.1447014, -0.0835920, 0.1993796, -0.2037404, 0.2378802, 0.0733893, 0.1031246, -0.1720252, -0.1576961, -0.1577295, 0.1765937, 0.1549924, 0.2782370, -0.1794447, 0.0118224, 0.0386235, 0.1686083, -0.0455125, 0.0239479, 0.3363706, 0.2048784, -0.1514463, -0.1784110, -0.0554486, 0.1295304, 0.0243738, -0.1712240, 0.2972542, 0.0428932, -0.0114672, -0.0491681, -0.0554807, 0.1232410, 0.0568912, 0.1307393, -0.2093795, -0.0658556, -0.0678602, 0.0588753, 0.2136323, 0.3961758, 0.2530802, 0.3053375, -0.2094321, -0.0534984, 0.3255486, 0.0317134, 0.2604698, -0.1292558, -0.2313743, 0.5022756, -0.1280835, -0.1903213, -0.1675902, -0.0633749, 0.2253595, -0.0438080, -0.0441033, 0.1290031, 0.0155377, 0.1203238, 0.0298378, -0.0318548, -0.1738139, 0.3517854, 0.2397738, -0.1761221, -0.0694951, -0.1605873, 0.2062358, -0.0374226, 0.1420348, 0.3723019, -0.0568254, -0.0438173, -0.1258350, -0.0595292, -0.1110766, 0.3408914, -0.2055839, 0.3553964, 0.3779454, 0.1820269, -0.3713968, -0.1388907, -0.0583377, -0.2509928, 0.3726457, -0.2565315, -0.2500832, 0.6859808, -0.0939390, -0.3671419, -0.1182951, -0.4170281, 0.3656015, -0.1447130, -0.3589243, 0.3429971, -0.3666881, -0.0388500, -0.1183596, -0.2116248, -0.1762650, 0.3876765, 0.1246309, -0.1588017, -0.1716887, -0.2300313, 0.5103440, -0.1204231, 0.3545428, 0.3863472, 0.1325386, 0.1332883, -0.0364773, 0.0036845, 0.0007496, -0.0258561, 0.1139374, 0.1049101, -0.0055429, 0.0586845, 0.1560625, 0.1160577, 0.1106960, -0.0156630, 0.0826044, 0.1043653, -0.0026794, 0.0908673, -0.0543923, -0.0376300, 0.0673608, -0.0336134, -0.0890906, 0.0366799, 0.0758745, 0.1865144, 0.0902447, 0.0911610, 0.2670291, 0.1246753, 0.0521441, -0.0851861, 0.0002922, -0.0310630, -0.1160178, 0.0275236, -0.0821817, -0.0199972, 0.0672117, -0.0605846, -0.0729758, 0.1130812, 0.1269108, 0.0561202, -0.0258951, 0.1678156, -0.0371948, -0.2252202, -0.0821187, -0.0521155, 0.1216106, 0.0768186, -0.2434731, -0.1177112, -0.2321903, 0.0542161, 0.0463736, 0.0254532, 0.0924203, 0.0517488, 0.1362362, 0.0411981, -0.0076017, 0.0303350, -0.0481525, -0.0132699, -0.0159446, 0.0674907, 0.1290068, -0.0090871, 0.0961170, 0.1847133, 0.0255950, 0.0076374, -0.0435950, 0.1342888, -0.0053795, 0.0688614, 0.1808659, 0.0809137, 0.0257069, 0.1353322, 0.0684837, 0.0528254, -0.0271843, -0.0789289, 0.2348697, -0.0137017, -0.0590185, -0.0944515, -0.0482381, 0.2542883, -0.0164956, -0.1154247, -0.5354905, -0.1545325, -0.0728251, 0.2142532, 0.0601069, 0.0387758, 0.0084679, -0.0490019, -0.2128936, 0.1065804, -0.0827505, 0.1655410, 0.0177874, 0.1086737, 0.2009658, -0.0532570, -0.0024164, 0.0842366, -0.1658569, -0.2513256, 0.0171698, 0.2903182, -0.0055659, 0.0502733, 0.0349598, 0.0711115, 0.1213169, 0.1131479, -0.5208188, 0.1984240, -0.0454542, -0.7446180, 0.2436450, 0.1842843, -0.1209646, 0.2367419, -0.0377841, -0.1012051, 0.1464775, 0.0640338, 0.1529063, 0.0851315, -0.0723902, 0.0897400, -0.0814293, 0.3493865, -0.2788113, 0.2167479, 0.0585168, 0.1732862, 0.4089991, -0.0716810, 0.4109166, 0.2199213, -0.0944595, 0.1484776, -0.0904212, -0.1657053, 0.0789018, 0.2197544, 0.1296805, -0.0744212, -0.3905227, 0.1584817, -0.5938300, 0.1462564, 0.0725910, 0.1132845, 0.1610459, -0.0708519, 0.0719044, -0.0301351, 0.2899398, -0.3059565, -0.0619260, -0.0280547, 0.1076971, 0.0561828, -0.1629360, 0.0200853, -0.2801204, -0.0455254, 0.0417354, 0.2537169, 0.0235625, 0.0960304, 0.0331727, 0.0438474, -0.0860837, 0.0537701, -0.0370125, 0.1101862, 0.1134432, 0.0725072, 0.0602296, -0.0669360, 0.0152163, 0.1004122, 0.0024781, -0.1365606, 0.0383805, 0.3197757, -0.0050766, -0.0110819, 0.0251403, 0.1252665, 0.0049781, 0.1642458, -0.4939194, 0.0236181, -0.2095826, -0.3558587, 0.3471970, 0.2901908, 0.2228802, 0.4416845, -0.4405195, -0.1233012, 0.2433387, 0.0972252, 0.2605558, -0.1425552, -0.3481513, 0.2001454, 0.0023520, 0.0956471, -0.5776583, 0.0427856, 0.2990909, 0.0509003, 0.2037649, -0.2108330, 0.1793235, 0.1205079, -0.3735260, -0.1639340, -0.3849420, 0.2819736, 0.2321640, -0.1131504, 0.2124343, -0.2218775, -0.0216871, -0.0267743, -0.2125342, 0.5066826, -0.0006396, 0.0969330, 0.0739221, 0.0080511, 0.0119026, 0.1029029, -0.0188758, -0.2749955, -0.0752128, -0.0558853, 0.0477102, 0.1539991, -0.1024775, -0.0638848, -0.1975829, 0.0218575, -0.0285837, 0.0232391, 0.0387695, -0.0237096, 0.1672437, -0.1230370, -0.1731672, 0.0753675, -0.2149828, 0.0464351, -0.0650896, 0.0355101, 0.1693525, 0.0077190, 0.0703532, 0.1099768, -0.2141089, -0.0487381, 0.0536241, 0.0519105, 0.0613161, 0.0489378, 0.1606165, -0.0225145, 0.0466986, -0.0501445, 0.0346053, 0.0145483, -0.0499784, 0.1480622, 0.0466610, 0.2586126, 0.1372464, -0.0182064, -0.0080250, 0.0357067, 0.1421851, -0.1336727, 0.2172560, -0.1339311, -0.1008614, 0.2790274, 0.0439150, -0.1276394, -0.1088914, -0.0811846, 0.1772669, -0.0211612, 0.0177003, 0.1642864, -0.1061374, 0.0523854, 0.1079330, 0.0232225, -0.1101582, 0.1603822, 0.0320467, 0.0091489, -0.0507098, -0.0115780, 0.1501948, -0.0699283, 0.1223872, 0.0706037, 0.1724578, 0.2006493, 0.0649078, 0.1509668, -0.0623790, -0.0645511, 0.1808354, 0.1149253, -0.1154514, -0.1008294, 0.1451701, -0.0502675, 0.0752371, -0.0804128, 0.0006339, 0.0477578, 0.0035055, 0.2220390, -0.0301222, -0.0329600, -0.0576776, -0.0689740, -0.2422004, 0.0937575, -0.0099750, 0.2292543, -0.0517892, 0.1508190, 0.1840941, 0.0448145, 0.0113271, -0.0087870, -0.2098651, -0.0405319, -0.0865703, 0.0608525, -0.1214489, 0.1369526, 0.0264936, -0.0173321, 0.2467832, 0.1529957, -0.1450258, 0.1439419, 0.0351723, -0.2249118, 0.2941892, 0.2552981, 0.0236458, 0.0462854, 0.2515261, -0.3204952, 0.2148926, -0.0329194, 0.2630965, 0.1989741, -0.0368212, 0.4208713, -0.3800537, 0.0155176, -0.0740606, 0.1267790, 0.0419056, 0.1632339, 0.1606868, 0.2138847, 0.1911425, 0.2951009, 0.1560645, 0.2185929, 0.0584907, -0.2082999, 0.0865987, 0.0716124, -0.3021580, 0.0203753, -0.2196450, 0.1195723, -0.0520162, -0.0265863, 0.0389293, 0.1018264, -0.0939442, -0.0325227, -0.1253860, -0.0749359, 0.0922435, 0.0995303, -0.0531026, -0.0457044, -0.0688948, 0.0230790, 0.0922221, -0.0824786, -0.0255360, -0.0129951, -0.0829752, 0.0937050, 0.0186503, -0.0806133, -0.1307621, -0.0972282, -0.0692211, 0.0582317, -0.0116887, 0.1092325, -0.1120776, 0.1327256, 0.0463738, -0.0787693, -0.0662544, 0.0855845, -0.1006780, -0.1527360, -0.0340169, -0.0687556, -0.0591476, -0.0022611, 0.0138223, 0.0629551, 0.1380066, -0.0126510, 0.0977846, 0.1045076, 0.0989738, 0.0377657, -0.0811700, 0.0202605, 0.0915152, -0.0039824, 0.0510247, -0.1335782, -0.1464067, -0.1585859, 0.1777178, 0.0189110, 0.0827761, 0.0979859, -0.0461295, -0.0075076, 0.0256631, -0.0288955, 0.0683214, 0.0877428, -0.0392019, 0.0710391, -0.0407132, -0.0602790, 0.0081490, 0.0073108, 0.1140437, 0.0012585, 0.0260943, 0.0574515, -0.0751549, -0.0177831, 0.0940683, 0.1106618, 0.0743542, 0.0056808, 0.0487135, 0.0444876, -0.0412027, -0.2176487, -0.0408573, 0.1326992, 0.1360583, 0.1574319, -0.0087728, 0.0350326, 0.0383005, 0.1677301, -0.0899560, 0.0603665, -0.0259673, -0.2500352, -0.0972897, 0.0987214, -0.0327828, -0.0035952, 0.1426999, -0.1058758, -0.1273733, 0.0268831, -0.2070621, 0.2052089, -0.0231421, 0.0271448, 0.2634265, 0.0220661, 0.0907134, 0.1305811, -0.0349100, -0.3506555, -0.0841024, 0.0707901, 0.0669807, -0.2059292, 0.1305924, -0.0017671, -0.1058832, 0.1278617, -0.1149769, -0.1362939, -0.1204103, -0.2196649, 0.2215740, 0.2071535, 0.2603668, 0.3312128, -0.3669798, -0.0984456, 0.2412032, 0.1198529, 0.1883393, -0.1618023, -0.1499168, 0.1292518, 0.0526435, 0.1848968, -0.4160731, -0.0300654, 0.2207760, -0.0654240, 0.1989535, -0.1675083, 0.2636143, 0.1874060, -0.3118060, -0.2380140, -0.1439105, 0.2592799, 0.2193761, -0.2358992, 0.1271154, -0.1230484, -0.0117411, -0.1407662, -0.0970296, 0.3945418, -0.0521388, 0.1640701, -0.0377531, 0.0156234, -0.1340219, 0.1431003, 0.2116156, -0.0530965, 0.0195240, 0.1177374, 0.0435956, 0.0355136, 0.0378757, 0.0067227, -0.0855447, -0.1282612, -0.0872343, 0.1607592, 0.1653295, 0.0517269, 0.0049176, 0.0341877, 0.0342692, 0.0820816, 0.2474246, 0.1051557, 0.1297041, 0.1552577, -0.0243321, 0.0605974, -0.0957303, 0.1119139, 0.0997945, -0.0398918, -0.0431664, 0.0971450, 0.1159252, -0.0556577, 0.0176815, 0.1574398, -0.0368445, 0.2868530, -0.1071068, 0.0065098, -0.3005257, 0.1361497, 0.1523075, 0.2592051, 0.1427121, 0.0577772, 0.1275293, -0.2132002, 0.1272033, -0.2412871, 0.1295094, 0.0751245, -0.1802343, 0.4050291, -0.1119642, -0.2620651, -0.2264495, -0.0372455, 0.1391363, 0.0483189, -0.0483137, 0.0681028, -0.1377683, 0.3082125, 0.1766223, -0.1050549, -0.2528051, 0.1726071, 0.2360788, -0.2281096, -0.3017775, 0.0190179, -0.0218340, 0.0789787, 0.1970388, 0.3049650, -0.0278723, 0.0756930, 0.1618495, 0.0722008, -0.0031999, 0.2081428, -0.0957281, -0.3623457, -0.0059590, -0.0567353, 0.0824867, 0.1861339, -0.2918355, -0.1380417, -0.1464277, 0.0028127, 0.0089564, 0.0760901, 0.0481130, -0.0057165, 0.2343063, -0.0907090, -0.1084133, 0.0491015, -0.2118946, -0.0320084, -0.1160605, 0.0060376, 0.1524979, -0.0489798, 0.0380263, 0.1805392, -0.0994991, -0.0714556, 0.0373607, 0.0946551, 0.1432712, 0.1358280, 0.1801252, -0.0144708, 0.0552264, -0.1420590, -0.0286320, 0.0409646, 0.0310048, 0.0688170, 0.2401502, 0.2150135, 0.1024110, 0.1378750, 0.0439814, -0.0845282, 0.0633488, 0.0049144, -0.0144915, -0.0112389, -0.0058419, 0.4445570, -0.2934993, 0.0578635, 0.0604731, 0.1893413, 0.1922132, -0.0107705, -0.1428461, 0.2218179, 0.2121445, -0.0839101, 0.0780201, 0.0436733, 0.0045098, 0.1067356, 0.1349622, -0.0093067, -0.1755681, 0.2301014, 0.0370817, -0.0517948, 0.1528491, 0.1649895, -0.1318644, 0.1311488, 0.0826844, 0.0368700, -0.1856733, 0.1061280, 0.0461970, 0.1590937, 0.1300075, -0.0080377, -0.0409849, 0.3044941, 0.0861371, -0.0561821, 0.0017463, -0.0597178, 0.0210516, 0.0111544, 0.1441629, 0.0214309, 0.0049699, -0.2185714, 0.0050840, -0.0408343, -0.0216587, -0.0164726, -0.1774084, 0.0590297, 0.0650206, -0.2016949, -0.0034298, 0.3638084, -0.0183775, -0.1294693, 0.0739247, 0.0509029, 0.1102410, 0.0299345, 0.0748930, 0.2274390, 0.0429069, 0.1959324, 0.0801827, 0.0925399, -0.0352699, 0.0183208, 0.1031433, 0.1881527, -0.1040827, 0.0212120, 0.1790782, -0.1017893, 0.1306964, 0.0237922, 0.1463627, 0.0948387, 0.0384656, 0.1718559, -0.0209177, 0.1101362, -0.0095538, 0.1117392, -0.0306590, 0.0564068, 0.0968896, 0.0729588, 0.0944791, 0.1225936, 0.1210719, 0.1033503, -0.0049769, 0.0287822, 0.0794007, 0.1234306, -0.0259578, 0.1317482, -0.0953752, 0.1388621, 0.0272338, 0.1188549, -0.0629802, 0.0412404, -0.0698351, -0.2295121, -0.1194893, 0.0438981, 0.1754096, 0.1712518, 0.0814118, 0.1364181, -0.1553219, 0.0363188, 0.1835890, 0.0181412, 0.0292746, -0.1994002, -0.1424536, 0.2042916, -0.0067361, -0.0845497, -0.1441885, -0.0365990, 0.0177396, -0.0433158, -0.0439082, 0.1204174, -0.0259898, 0.1197867, -0.1547542, -0.1143212, -0.0759045, 0.2180412, 0.1017659, -0.3494031, -0.0166721, 0.0119040, 0.1696634, -0.1999388, 0.0120715, 0.2797334, -0.0194539, -0.1313359, -0.0544571, 0.1231139, -0.0004430, 0.0079620, 0.0202534, 0.1094951, 0.1640913, 0.1317416, -0.0980887, -0.1546040, -0.0686703, -0.1390513, 0.1254304, -0.0875308, -0.0082511, 0.1624585, -0.0752121, -0.0355348, -0.1163182, 0.0141144, 0.1648181, 0.2056155, 0.1264143, -0.0289152, -0.0225983, -0.0597615, -0.1753401, -0.0436264, -0.1789621, -0.0370500, 0.0757054, 0.1939042, 0.1418326, -0.0479703, 0.1574003, 0.1600773, -0.0139411, 0.0913531, 0.0098097, -0.1352293, -0.0796148, -0.1194437, 0.0490133, 0.0815637, 0.0929295, 0.1606549, 0.1790670, 0.1203449, -0.0485154, 0.0798035, -0.1198460, 0.1152097, 0.0411213, -0.2034393, -0.0118019, 0.1814440, -0.2090694, -0.0012390, 0.0934856, 0.0496952, 0.1510418, -0.1059456, -0.2545933, 0.1221723, 0.1059813, -0.1581935, -0.0107117, 0.0093857, -0.0051760, 0.1763689, 0.0836858, -0.1396340, -0.1494944, -0.0327679, 0.1106670, -0.1474925, 0.1469030, 0.1235508, -0.0984524, 0.1817849, 0.0194061, -0.1091003, -0.3327752, 0.1195140, 0.0988613, 0.1214290, -0.0291529, 0.0945024, 0.1112337, -0.0306930, 0.0743293, -0.1953720, 0.1601515, 0.1445819, -0.0352879, 0.1118519, -0.0652564, 0.0496083, -0.0637741, -0.0705349, 0.0367163, -0.0375448, -0.0140134, -0.0080775, -0.0903875, 0.2063550, 0.1241419, -0.1003668, 0.0145737, 0.0811796, 0.1637033, -0.1318309, -0.2958232, 0.1483957, -0.2284489, -0.1507302, 0.1874386, 0.1962604, 0.1345763, 0.0032363, 0.1621924, 0.3156036, 0.0221805, -0.1051835, 0.1644241, -0.0268363, 0.0951453, -0.1128005, -0.0587732, 0.1955625, -0.0377200, -0.1108181, -0.0957728, -0.3910260, 0.0068945, 0.2859435, 0.0915639, -0.1549890, -0.0977180, 0.1199048, 0.1356267, 0.2200986, -0.0310339, 0.0940667, 0.0140953, -0.0184307, 0.1553808, -0.1161039, -0.3301682, 0.2545203, -0.0440544, 0.0315271, 0.2519795, 0.1310226, 0.2259545, 0.3054750, -0.1189765, 0.1986749, 0.0344283, 0.0140387, 0.0703262, -0.0399852, 0.0595102, 0.0438197, 0.0557346, -0.0020117, 0.0873360, 0.0236786, -0.0484008, 0.1152349, -0.0569095, -0.0750718, -0.0206955, -0.0409074, 0.0643409, 0.1044797, -0.0196116, 0.0698416, 0.0684118, 0.0021101, 0.0889270, -0.0188106, -0.1380123, 0.0239174, -0.0255226, 0.0230307, 0.0038029, -0.0656509, 0.0443848, 0.0794129, 0.0412097, -0.0774947, 0.0314676, 0.1333432, 0.0383199, -0.0336161, 0.0806065, 0.1471461, 0.1621533, -0.1251352, -0.0131962, 0.0210453, 0.1548973, 0.0537133, 0.0223532, -0.1264131, 0.1144637, 0.1564578, 0.0815183, -0.0981182, 0.0133031, 0.0863826, 0.1981653, 0.0547608, 0.0473645, 0.0773910, -0.1341602, 0.0623165, 0.0924456, 0.1088680, 0.0257381, 0.0160282, 0.0596595, 0.0189063, 0.1636666, -0.1186088, -0.0421625, 0.1842708, 0.1642664, -0.1521130, 0.1478984, 0.0601312, -0.0989925, 0.0400505, -0.0538377, 0.0098670, 0.0294296, -0.1165547, 0.1754065, -0.4778605, -0.2941010, 0.1447939, 0.2513632, -0.0188511, 0.0823858, -0.2938265, 0.0505118, 0.2602015, 0.2345427, -0.1180933, -0.1884277, 0.3315710, 0.2555118, 0.1797279, 0.1327202, 0.0653798, -0.3106444, 0.1991696, 0.2355832, 0.2427837, 0.1746736, 0.1483534, 0.3142463, 0.1180298, 0.3673099, -0.4951557, 0.0793610, 0.6057323, 0.2512293, -0.3050209, 0.2356037, 0.3647200, -0.1129147, -0.0218021, -0.1453494, 0.1170148, -0.1163395, -0.1813274, -0.0261384, 0.1960459, -0.0274579, -0.2188147, -0.0563061, 0.2414129, -0.1184785, 0.1718882, 0.1935556, 0.0126834, 0.1518441, 0.2302544, 0.1066893, 0.1098915, 0.1130985, 0.0986460, -0.0247016, 0.0928637, 0.2377490, -0.1032502, 0.2000188, -0.0812773, -0.0289391, -0.1874364, -0.0280817, 0.2900079, -0.0535570, 0.2057519, 0.0539481, -0.1427161, 0.0067021, 0.3520680, 0.1103427, -0.0876207, -0.0968005, -0.0423117, 0.0930265, -0.1996089, 0.1001825, 0.1617280, -0.0969321, 0.2663080, 0.0925281, 0.0106847, -0.1795804, 0.1949377, 0.0131001, 0.1614010, -0.0324339, -0.0775544, 0.0828635, 0.3230765, -0.0119157, -0.0302509, -0.1076361, -0.0883691, -0.0133969, 0.0276654, 0.2711909, -0.0352767, 0.0777718, -0.0885241, -0.0764456, -0.0107692, -0.0271117, -0.0019054, -0.1276367, 0.1076251, 0.1696165, -0.1402323, -0.1251156, 0.4237353, -0.0645978, -0.1446269, 0.0562831, 0.2159663, 0.0391100, 0.0033314, 0.1322868, 0.1872354, -0.2398212, 0.3096692, -0.0175039, 0.2847298, -0.3441766, 0.1796474, 0.1290699, 0.1575038, 0.0107287, -0.0026415, 0.0551120, 0.0051556, 0.1590871, -0.2930738, -0.1323932, -0.1056955, -0.1023347, 0.3105602, 0.1812643, -0.1373847, -0.2132123, -0.0421029, 0.1634240, 0.1659188, 0.0843617, 0.1735548, -0.1633014, 0.1823196, 0.0454075, -0.0627089, -0.2283692, 0.2882977, 0.1162156, -0.0264279, -0.0157533, 0.1066637, 0.1250917, 0.3921202, 0.0853172, 0.3117524, -0.2983531, 0.0962090, -0.1266262, 0.2786442, -0.2460207, 0.0736843, 0.0303346, -0.0958560, -0.0365098, 0.0476499, -0.0533397, -0.0845239, 0.0185575, 0.0021276, -0.0249386, -0.1315887, -0.1158995, -0.0291226, 0.1372428, 0.0054620, -0.2074444, -0.0137355, 0.1331849, 0.4169787, 0.5479227, -0.2323936, -0.0303335, 0.0048643, -0.1707017, 0.0184426, -0.2963170, 0.1182924, 0.1411022, 0.2567138, 0.4380273, -0.1468389, 0.1372215, 0.2733213, -0.2153721, 0.2453651, 0.1169594, -0.6139002, -0.1810029, 0.2275981, 0.1928892, -0.2921035, 0.2601596, -0.3773378, 0.1329535, 0.1126974, -0.0190404, -0.0407438, -0.1037840, 0.2279289, 0.0705745, 0.0059767, 0.1146948, 0.2375422, -0.3720233, 0.0330309, -0.0247462, 0.1263302, 0.0855027, 0.1514393, 0.2401773, 0.1511949, 0.2466107, -0.4319224, -0.0314389, 0.3353460, 0.1272511, -0.3015556, 0.0700754, 0.2389252, -0.1266733, -0.0341708, -0.1185521, 0.1635069, -0.1181192, -0.0147705, -0.2589327, -0.0535843, -0.0678646, -0.0292926, 0.0150273, 0.2309411, -0.2090789, 0.0700409, 0.1216534, 0.2626362, 0.1477809, 0.0984420, -0.0513403, 0.2248360, 0.2150395, 0.1588731, 0.0636056, -0.1531290, 0.0373994, 0.2667404, 0.1649891, 0.0225995, 0.2026966, -0.1494437, 0.0220558, -0.3598399, 0.1083493, -0.0640293, -0.1713031, 0.1628814, 0.1613757, -0.0999689, 0.2621071, 0.1720401, -0.0811750, -0.0667860, -0.0435994, -0.0817527, 0.0545733, -0.0663439, 0.1746157, -0.0614617, 0.0421815, -0.0267600, 0.2573066, -0.2179244, 0.1334192, -0.3336070, 0.1924198, 0.1175023, -0.1405872, 0.1049479, -0.1024917, 0.2348744, 0.1062307, -0.0866145, 0.0958758, 0.1482157, -0.0407248, 0.0612788, 0.0417245, 0.0367123, 0.0940546, 0.0747358, 0.0170333, -0.0068363, 0.1207409, 0.0288141, -0.1097021, 0.0376890, 0.0753941, 0.0175572, -0.0958828, 0.0390824, 0.2038161, 0.0093829, 0.1071602, 0.0042600, 0.0287114, 0.0943354, 0.1390502, 0.0020709, 0.0575044, -0.1062860, 0.0915635, -0.0414735, -0.0002831, 0.0408632, 0.0397658, 0.0702590, -0.1584304, 0.0247971, -0.0131415, 0.0726104, 0.0500959, -0.0192518, 0.0250406, 0.1171361, -0.0394304, -0.0201220, -0.0006755, -0.0935123, 0.0089302, -0.0389297, -0.2013032, 0.0395240, -0.0066659, 0.0377690, -0.0767429, -0.0223380, 0.0607305, -0.0140283, -0.0546392, -0.1016295, 0.0647305, 0.0219167, 0.0489217, -0.0489016, 0.0520324, 0.0492256, -0.6348464, 0.0266418, -0.3675595, 0.0430778, -0.3648075, 0.2725258, -0.0338469, -0.3297566, 0.0129249, 0.1551451, 0.1829595, 0.0749601, 0.0780471, 0.2387420, -0.1716642, -0.1171492, -0.1202646, -0.1162516, 0.1647016, 0.1093555, 0.0406478, 0.1285902, 0.1717578, 0.1942453, 0.8117667, -0.4531624, 0.1020376, -0.0212048, -0.0545113, 0.0752259, -0.3427546, 0.0944520, 0.2675176, 0.1158641, 0.3697310, -0.1470877, 0.1957724, 0.1043548, -0.5287858, 0.1211028, -0.1874333, -0.1272655, -0.1321331, 0.1594464, 0.0120122, 0.0895118, -0.1230484, -0.3218101, 0.0554665, 0.1254307, 0.2292020, -0.1707701, -0.1685847, 0.0814393, 0.0785623, 0.1957546, 0.1095330, -0.1574423, -0.1101131, 0.2359957, 0.1256229, 0.1786378, 0.1558309, 0.1014782, 0.2494805, -0.0196141, 0.1911481, -0.1970124, -0.0381590, 0.3419618, 0.0913707, -0.2050981, 0.2366614, 0.4030797, -0.2272097, -0.0250007, -0.1912125, 0.1842245, -0.1653676, -0.1163872, -0.2053791, 0.3309465, 0.0791354, -0.1666836, -0.0090151, 0.4439151, -0.4528796, 0.0780491, 0.0125575, 0.1430468, 0.1162437, 0.1390403, 0.0001863, 0.0963567, 0.2475069, 0.4114440, 0.0683822, -0.3577030, 0.3374866, 0.2151009, 0.4038861, -0.1049911, 0.1417068, -0.2987642, 0.1617424, -0.1935217, -0.0071909, 0.0719540, -0.2155504, 0.0373235, 0.4342237, 0.1013507, 0.2509070, 0.1620697, -0.1496994, -0.1249816, -0.2397861, -0.2320750, 0.3162317, -0.0332510, 0.0048704, -0.0863008, -0.0092617, -0.0667787, 0.0022336, 0.3105580, -0.0114588, 0.4372088, 0.1242324, 0.2341002, 0.0558579, 0.0676831, -0.0432284, -0.0450027, 0.2733792, 0.0484995, -0.0331210, 0.2542304, -0.0111942, -0.1023124, 0.1064168, -0.0595995, 0.1892952, -0.0599754, -0.0433932, 0.3131855, -0.0542501, 0.0076646, -0.0429329, 0.0253939, -0.1285302, 0.3530476, 0.1814922, 0.0329953, 0.0550926, -0.1153610, 0.1413730, 0.0372003, 0.2079058, 0.2171673, -0.4153239, 0.0998747, 0.2256052, 0.4492763, -0.4389136, 0.2717132, 0.1277074, -0.0590417, -0.1238914, 0.0130654, -0.0454077, -0.1558806, -0.1029910, -0.4871519, -0.2158463, -0.2391966, -0.1357863, 0.3264276, 0.1760900, 0.0570249, -0.3804869, 0.0741366, 0.3852479, 0.4246385, 0.3162591, -0.3173400, -0.1612527, 0.1517522, -0.0887173, -0.1303628, -0.2834306, 0.2331056, 0.2961074, 0.1054189, 0.2030887, 0.4475395, -0.0388273, 0.6836708, 0.2229970, 0.5330814, -0.4718321, 0.0197487, -0.2296067, 0.3489790, -0.3781360, 0.2112288, -0.0449259, -0.1746838, -0.3095363, 0.0452265, 0.0465521, -0.1168272, -0.0513902, -0.2699390, -0.1903950, -0.0515170, -0.2229921, -0.0027608, 0.1463737, 0.1177083, -0.1006469, 0.1689691, 0.0828116, 0.4010498, 0.5519857, -0.3771348, -0.0428920, -0.0555358, -0.1412400, 0.2475460, -0.2190264, -0.0321716, 0.1312060, 0.4117754, 0.2716603, 0.1398298, -0.0425524, 0.3154992, -0.2185508, 0.1964961, -0.0789269, -0.1583173, -0.1351647, 0.2750350, 0.0315003, -0.1846549, 0.0347652, -0.5048093, -0.1312642, 0.0812051, -0.0074290, -0.1118369, -0.1686248, -0.0004670, -0.0591206, 0.0972121, -0.0172256, -0.0682763, -0.0281533, 0.1802052, 0.0183115, 0.1345306, 0.0156171, 0.2045158, 0.3553780, -0.0987021, 0.1107653, -0.1728431, -0.0173259, 0.3679817, 0.0962263, -0.2991435, 0.0888769, 0.2963883, -0.1334020, -0.0173164, -0.2481795, 0.2876331, -0.1089204, 0.0425519, -0.3402748, 0.1117289, -0.1121095, -0.0179950, -0.0341042, 0.0940629, -0.2576209, 0.0116677, 0.1206662, 0.1636565, 0.0433948, -0.0812420, 0.0686592, 0.0875186, 0.3295775, 0.1761509, 0.0407536, -0.1160521, 0.0631372, 0.0573396, 0.0415582, -0.0465808, 0.2798915, -0.0844449, 0.1168608, -0.5493878, -0.1330620, -0.0073455, -0.2525773, -0.0761991, 0.1389131, -0.1458222, 0.1905272, 0.1543743, -0.0314543, -0.2375194, 0.0577378, 0.0454281, 0.0840030, -0.0124640, -0.0657277, 0.1361820, -0.1228325, 0.0696939, 0.0070158, -0.0516439, 0.1132289, -0.4117408, -0.1130808, 0.0703485, 0.0981867, 0.1260078, -0.0119312, 0.1602790, -0.1299283, 0.0772723, 0.0090652, -0.1202663, 0.2208068, 0.0908430, 0.0124919, 0.0500531, 0.0571967, 0.2673512, 0.2917509, -0.1023982, 0.2445126, 0.0532292, 0.0837670, 0.2119151, 0.0757254, 0.0728718, -0.0549590, 0.1405547, 0.2308909, -0.0580344, -0.0134771, 0.1528948, -0.1682475, 0.0407296, 0.0535979, -0.1461451, -0.0399139, 0.0490499, 0.0601362, 0.0196799, -0.0962559, 0.1542039, 0.1636334, 0.1192503, -0.1411506, -0.0858464, -0.1478281, 0.0296560, 0.1563600, 0.0452051, 0.0347293, 0.1452560, -0.1118490, -0.0213240, -0.0140103, -0.0448858, 0.1728302, -0.0064842, -0.1921436, 0.0603268, 0.0268588, -0.0465377, -0.0983047, 0.0864975, 0.1095269, -0.0140637, 0.1058367, 0.0788052, 0.0257851, -0.2032152, 0.0591213, 0.0966469, 0.0571464, -0.0157513, -0.5763256, 0.1383430, -0.3985586, 0.1394826, -0.4277131, 0.2202266, 0.0757168, -0.2274538, -0.1343325, 0.1106775, 0.1178819, 0.0203526, 0.2212098, -0.0467066, -0.2167545, -0.1436238, -0.3252617, -0.1022794, 0.1991487, 0.0482763, -0.0074843, 0.0790763, 0.1676632, 0.4736833, 0.9084331, -0.4185829, 0.0613974, 0.0041251, 0.0466121, -0.0529079, -0.4578123, 0.1078048, 0.2343530, 0.1566904, 0.6802756, -0.1426113, 0.1697837, 0.2171997, -0.4484621, 0.1781316, 0.1942663, 0.0007670, -0.0096135, 0.0437983, 0.1018373, -0.0926703, 0.1463403, -0.0732209, 0.0122584, -0.0557905, 0.0776975, 0.1069728, 0.0134866, 0.0843047, -0.0070934, 0.0473517, 0.0636259, 0.0564047, -0.0985624, 0.0714485, 0.1859832, -0.0245172, -0.0183365, 0.1387494, 0.0110663, 0.1129785, 0.1936160, -0.0616369, 0.2242678, 0.1133951, 0.0624081, -0.0949640, -0.0210500, 0.0436100, 0.0185977, 0.1043095, -0.0280889, 0.0416746, 0.0182676, -0.1233193, -0.1173006, 0.1640717, 0.0244871, -0.0753799, -0.0220871, 0.0696501, -0.0029220, 0.0175979, -0.1534093, -0.0057806, -0.0454661, -0.0361456, -0.0207257, -0.0308917, -0.0065107, 0.0902464, -0.0353312, -0.0180289, 0.1468765, 0.0681654, -0.0575691, -0.1201942, -0.0428579, 0.0406337, -0.1010535, -0.0826630, -0.0458272, 0.1793382, -0.0111534, 0.0231708, 0.0913504, -0.0006291, 0.0058579, 0.0003548, 0.0575857, -0.0494074, -0.0994353, 0.0221827, 0.1130704, 0.0776482, 0.2729671, -0.1827839, 0.0840648, 0.0739232, 0.1422416, 0.0471722, 0.2660519, -0.0095864, 0.1609224, 0.2097572, 0.3070095, 0.0784734, -0.0193643, 0.1797003, 0.1229597, 0.2048974, 0.1240609, 0.1482985, -0.2165084, 0.1478706, 0.3064558, 0.2338981, 0.1232074, 0.1707039, 0.2445283, 0.2218673, 0.2739997, -0.1677472, 0.1270156, 0.2494890, 0.0577390, -0.0174810, 0.2135214, 0.1675759, -0.1272914, 0.1464084, 0.0063575, 0.1107919, 0.0756356, -0.0914719, -0.0457282, -0.0194779, -0.0835161, 0.1993377, -0.0899289, 0.0942539, 0.1040589, 0.0589800, -0.0077981, 0.1658010, 0.1099775, 0.0454760, -0.0056729, -0.0019395, -0.0741365, -0.0264836, -0.1672933, 0.1543074, 0.1639804, 0.0387975, 0.0837714, 0.1090338, 0.0220363, 0.1569429, 0.2224266, 0.0157026, 0.0932197, -0.0740852, 0.1788915, 0.1890251, -0.0574672, 0.1816876, 0.1024420, 0.1593503, 0.2493743, 0.1848412, 0.1037864, 0.1617894, 0.0190005, 0.1080146, 0.0518385, -0.0541828, -0.0403827, 0.0927396, 0.0364579, -0.0388541, 0.2050390, 0.0549149, -0.0061914, 0.1264973, 0.0228511, -0.1089097, 0.0432970, -0.0155725, -0.0103915, 0.0506506, -0.0333644, 0.2553892, -0.0436555, 0.0865601, 0.0535058, 0.0245737, 0.1058862, 0.1652154, 0.1058937, 0.1769238, 0.1276584, -0.0445110, 0.1770644, 0.1155222, 0.0493589, -0.0739788, 0.0633063, 0.0568524, -0.0428580, 0.0393320, 0.0010848, 0.0928586, 0.1333491, 0.0803015, -0.0707715, 0.0513050, -0.0350852, 0.1437939, -0.0219114, -0.0608836, 0.0236845, -0.0748551, -0.1297910, -0.2152590, 0.1298485, 0.0879284, 0.0392115, 0.0669349, -0.1120410, 0.0875246, -0.0412681, -0.1577983, 0.0538869, -0.0568869, 0.0627464, -0.0237062, -0.1608486, 0.1552377, 0.1241201, 0.0015989, -0.0997543, 0.1021652, 0.2170620, 0.1244571, 0.0233833, 0.0145548, -0.1057611, 0.1549796, -0.0271375, -0.0558862, 0.0064236, 0.1102640, -0.0954083, -0.1904996, 0.0500016, -0.0604231, -0.1406970, -0.0632834, 0.0154675, 0.1960555, -0.0400278, 0.0596844, 0.1482634, 0.3597887, 0.0112013, -0.2167898, -0.0580288, -0.0019081, 0.1706668, 0.0632613, 0.0448282, 0.0678205, -0.1768706, 0.1337608, -0.0156998, 0.1314189, 0.2346841, -0.0080859, 0.0552897, -0.1568744, 0.1708738, 0.0001708, -0.2393998, 0.1380935, 0.1167944, -0.0846671, 0.2749509, 0.0620462, -0.0457919, 0.0232058, -0.0097432, -0.0009463, 0.0183997, 0.1470320, -0.0152312, -0.0127884, 0.0024958, 0.0115063, 0.0368619, -0.0559453, -0.0638221, -0.0848354, -0.0702744, -0.2326523, 0.0757468, 0.0626536, 0.0325143, 0.0663108, -0.1062662, 0.0617895, 0.0929575, -0.0280942, 0.0237540, -0.0719248, 0.1211969, -0.1226605, -0.1831507, 0.0301497, -0.0098846, 0.0837976, -0.1548435, 0.0541723, 0.2229033, 0.1035980, 0.0981579, -0.0429075, -0.1683482, -0.0041653, -0.0439871, -0.1734778, 0.0190906, 0.0912377, -0.0367416, -0.2282218, 0.1182251, 0.1492234, -0.0068935, 0.0934384, 0.0137759, 0.0022735, 0.1545867, 0.1110216, -0.0437226, -0.0342445, 0.0868572, 0.1820915, 0.0960988, 0.1366398, 0.0617184, 0.1047327, 0.1461563, -0.0115561, 0.0989558, 0.1674807, -0.0459882, 0.0786214, 0.0322925, 0.1147922, 0.2487893, -0.0203824, 0.1444111, 0.1928886, 0.0313462, 0.0969312, 0.0557484, 0.0437703, 0.0022596, 0.1342676, 0.0410409, 0.0008705, -0.2161846, 0.0484170, -0.0343859, 0.1620306, 0.0181391, -0.1981987, -0.0545324, 0.0098197, -0.0229529, -0.0007966, 0.0468367, -0.0066748, 0.0167624, 0.0355006, 0.0115327, -0.1605519, -0.0536908, -0.0063705, 0.0179266, 0.0102955, -0.0584860, 0.0903738, -0.3086953, -0.0276340, 0.0207349, 0.0439633, 0.0252040, 0.0165736, -0.0205206, 0.0707061, 0.0975459, -0.1773454, 0.0410653, 0.0638787, -0.0218228, -0.0723969, 0.0111305, -0.0014910, -0.1064771, 0.0533918, -0.0028360, -0.0458553, 0.0380137, -0.0652859, 0.1481767, -0.0252765, 0.0557305, 0.0049973, 0.0511992, -0.0741908, 0.2029507, -0.2799301, -0.0471971, -0.1671384, 0.1765945, 0.2511335, -0.0523979, 0.1054301, -0.1760353, 0.0403918, 0.0549191, 0.0889212, 0.0383173, -0.0159798, 0.2159634, 0.0081386, -0.1951359, 0.1144471, 0.1419614, 0.2316262, 0.0517565, -0.1134935, 0.3958406, 0.0940323, 0.0312780, 0.0596914, -0.0866767, -0.0335487, -0.1077293, 0.0767812, -0.0271585, -0.0449044, 0.0007637, -0.1795420, -0.0560686, 0.1178853, -0.0892722, 0.0549485, -0.0370630, 0.0547381, 0.0582824, 0.0681430, 0.0238182, 0.2030651, 0.0286094, 0.0360454, 0.0122944, 0.1966252, 0.0589634, 0.1649318, 0.0264608, 0.0230437, 0.1743028, 0.0379246, 0.0623187, 0.0691725, 0.0623535, 0.0084008, 0.1260756, -0.1550827, -0.0102505, 0.1080355, 0.0362581, 0.1881656, 0.0776874, 0.2853732, 0.0814181, 0.0287903, 0.0160097, -0.1187789, 0.0201489, 0.0617338, -0.1112706, 0.2016945, 0.3034810, -0.0734822, -0.0672514, 0.1014831, 0.4208584, 0.0117990, 0.1952744, 0.1250204, 0.1631848, 0.4805285, 0.3695264, -0.2215645, -0.0025830, 0.2811304, 0.4870097, 0.5037735, 0.2625540, 0.1905249, -0.0987222, 0.3240893, 0.2880163, 0.5009637, 0.3694475, 0.0824161, 0.4379171, 0.0864480, 0.5036779, -0.0295229, -0.0168853, 0.4395336, 0.2969354, -0.1321647, 0.4847436, 0.4968588, -0.0510598, 0.0516762, -0.0419370, 0.0295255, -0.0229389, 0.0553524, -0.0822068, -0.0217808, 0.0404933, 0.0554144, -0.1245284, -0.0296280, 0.0635190, -0.0071062, -0.1374752, -0.1094643, 0.0252451, -0.0825683, -0.0169636, -0.1577899, -0.1646090, -0.0826430, -0.0567609, -0.0262780, 0.0017434, -0.0311532, 0.0065403, 0.0865867, -0.0442216, 0.0931917, 0.0536045, -0.2130326, -0.0507314, -0.0159146, 0.0091546, 0.0597620, -0.1060760, 0.0207395, 0.0171125, 0.0470834, 0.0605037, 0.1237045, -0.0495046, 0.1055468, -0.0939548, -0.0191632, 0.0386021, -0.0867955, 0.0059512, 0.0322966, -0.0058433, 0.0199676, 0.0648799, -0.0164399, -0.0051699, -0.0330469, -0.0197386, -0.0452983, -0.0744225, -0.0540695, -0.0318233, -0.0510204, -0.0492128, 0.0582954, -0.1260795, -0.0173263, -0.0179158, 0.0175982, -0.0142120, 0.0039859, -0.0266246, 0.0910552, -0.0179801, -0.1374286, 0.0802765, 0.0113738, -0.0165478, -0.0070872, -0.0040734, -0.0477625, -0.0853150, 0.0635534, -0.0042820, -0.0021926, 0.0160917, 0.0115308, -0.0543043, 0.0601115, -0.0206936, 0.0831114, -0.1053214, -0.0712914, 0.1889500, -0.1230636, -0.2249007, -0.1616038, 0.0056263, 0.2895736, 0.0582322, 0.0070477, -0.5623448, -0.0623202, -0.1169363, -0.0586280, 0.0873033, -0.0237504, 0.1181912, -0.0787659, -0.5570140, 0.1958815, 0.0587150, 0.2553654, -0.0312136, 0.0786364, 0.3256859, 0.0775414, 0.0199649, 0.1323861, -0.2384659, -0.0979230, 0.0267309, 0.0916445, -0.0190014, 0.0967229, 0.0330331, -0.1022071, -0.0504669, 0.0276000, -0.1678248, 0.2186421, 0.0110315, 0.1673816, -0.1025666, 0.1489910, 0.1533652, 0.3265910, 0.1676894, -0.2432321, 0.0581613, -0.0023584, 0.2071984, 0.1395652, 0.1128964, 0.0219564, -0.0528506, 0.2338562, 0.0715749, 0.2214495, 0.3044498, 0.0512893, 0.3233253, -0.2438018, 0.1864458, 0.0510733, -0.2275820, 0.2523723, 0.0943459, -0.1438199, 0.3901894, 0.3324445, -0.0053232, -0.0654641, -0.0883869, 0.1822854, -0.0677738, 0.1555850, 0.0821863, 0.0580648, 0.1205914, -0.1467984, 0.0714697, 0.0456437, 0.2087419, -0.2803899, -0.1301422, -0.2039494, 0.0903335, 0.3495255, -0.0029557, 0.1419024, -0.4152925, -0.0106836, 0.0044084, 0.0324887, 0.1475350, -0.0647783, 0.2780113, -0.1422167, -0.5672835, 0.1210460, -0.1033593, 0.2767604, -0.0493114, -0.0072320, 0.5451951, 0.0060682, 0.0564792, 0.0505406, -0.4343016, -0.2329224, -0.0033945, 0.1743140, 0.0768077, -0.0438748, 0.0267697, -0.2144765, 0.0316675, 0.2943739, 0.1183204, -0.0264360, -0.0118433, -0.0289546, 0.1755231, 0.1609333, -0.3143106, -0.0574546, 0.0654408, 0.3369988, 0.1423303, 0.0389881, -0.1506529, 0.0300340, 0.1644032, -0.1389041, 0.3113087, 0.3027665, -0.0657110, 0.0165073, -0.1877100, 0.1508706, 0.1586965, -0.0501889, -0.0246797, 0.2048583, 0.0053834, -0.0511851, -0.0442327, 0.3479496, -0.1189596, 0.0063904, 0.2662901, -0.0319677, -0.2265345, 0.1060596, -0.0908497, 0.2960060, 0.0330500, -0.2380487, -0.0015654, -0.0140934, -0.0028386, -0.0022547, -0.0319232, -0.0449213, 0.0133018, -0.0012581, 0.0010676, -0.1377882, -0.1043240, -0.0176294, -0.0132417, -0.0111195, 0.0000390, 0.0511653, -0.2216948, -0.0154148, 0.0081920, 0.0305609, 0.0049948, -0.0501286, -0.0201327, 0.0302302, 0.0383943, -0.2175659, -0.0198512, -0.0064076, -0.0007738, -0.0681973, 0.0420643, 0.0101024, -0.0623101, 0.0076651, -0.0224694, -0.0569942, -0.0021938, -0.0651182, 0.0931462, 0.0814887, 0.0542250, -0.0430116, -0.0632076, -0.0035832, 0.2770362, -0.0053792, -0.0733415, -0.0890590, 0.1622701, 0.3690603, 0.1085156, 0.0830341, -0.3429156, -0.0954893, -0.0674352, 0.1622930, 0.1848171, 0.0226873, 0.1623740, -0.0753543, -0.4376448, 0.1714128, 0.0550050, 0.2379043, 0.0086605, -0.0268659, 0.4615716, 0.0098489, 0.0024644, 0.2129045, -0.1798657, -0.2892630, -0.0189245, 0.1484560, -0.0058625, -0.0288026, 0.0528125, -0.0730481, 0.1774886, 0.1209675, -0.1344019, 0.2346229, -0.1249650, -0.0111982, 0.1849909, 0.2283492, -0.0696371, 0.0189871, 0.2862174, 0.0445547, 0.2061664, 0.1321106, 0.1765220, 0.1934761, -0.0272838, 0.2185779, 0.0436695, -0.0657933, 0.0378078, -0.0281314, -0.0949853, 0.2891657, 0.3819138, 0.1494023, 0.0264964, 0.1524735, 0.2630303, 0.3284010, 0.0171386, -0.0492094, -0.0025521, 0.1323384, 0.0105772, -0.2943521, 0.0216879, 0.2299275, -0.1842539, -0.0921848, 0.1757602, 0.3518650, -0.1850295, 0.1961615, -0.2090254, 0.0965816, 0.0433631, 0.4563712, -0.1366791, -0.0782589, 0.3109311, -0.0967063, 0.3675275, -0.0575650, 0.3526825, 0.3376830, -0.0877437, 0.4197026, -0.0788839, -0.2281028, -0.0441222, -0.2531815, -0.2143884, 0.2759043, 0.3004833, 0.0244051, -0.0915674, 0.2865615, 0.4816151, 0.2243564, 0.0709068, -0.0052964, -0.0094066, -0.0641138, -0.2715736, -0.1665811, -0.0661202, 0.1972277, -0.0569640, -0.0020929, -0.0544939, 0.1073532, 0.1329935, 0.1072376, -0.1560321, 0.0486212, 0.0482765, 0.0061501, -0.1860697, -0.0951641, -0.0090699, 0.0464260, 0.0355029, -0.0307318, -0.0437918, -0.0331203, -0.0120283, -0.0277294, 0.0810355, 0.0385793, -0.0199180, -0.1196606, -0.1080195, 0.1413427, -0.0149730, -0.0359332, -0.0844701, 0.0619313, 0.0397057, -0.0985200, -0.0392854, 0.0395540, -0.1697544, 0.0137045, 0.1072413, 0.0478157, 0.0432308, 0.0949292, 0.0209714, 0.0816406, 0.0691198, -0.3803334, -0.0615847, -0.0099157, 0.0428025, 0.0301442, -0.0157038, -0.0000884, 0.0500405, 0.0814076, -0.0381605, -0.0947569, -0.1153938, 0.0327580, 0.0437513, -0.0365241, 0.0057230, 0.0943574, -0.3829435, -0.0125963, 0.0406953, 0.0398517, 0.0787487, -0.0510762, -0.0295365, -0.0154967, 0.0602321, -0.2961187, -0.0352264, 0.0098716, 0.0359812, -0.0099290, 0.0632396, 0.0172901, -0.0596056, 0.0009392, 0.0006695, -0.0579372, 0.0087541, -0.0471119, 0.0739934, 0.0244656, 0.0961506, -0.0328566, 0.0261472, 0.0186900, 0.2029377, -0.2031569, -0.1091222, -0.0336411, 0.0005637, 0.1612643, -0.0956765, -0.0830001, -0.4552317, -0.0847095, -0.0738072, 0.0924278, -0.0717062, 0.0558137, 0.1895352, 0.0201376, -0.3046583, 0.0879356, -0.1539260, 0.2238764, 0.0545576, 0.0174300, 0.3519593, 0.0135685, 0.0570460, 0.0745141, -0.1494939, -0.1973537, 0.0309715, 0.3066823, -0.0248001, -0.0242831, 0.1639295, -0.0276248, -0.0921747, 0.2673063, -0.0313629, 0.1762896, -0.1611436, -0.1051114, 0.0678697, 0.0877446, -0.4854032, 0.0223404, 0.0791349, 0.0182178, 0.1418231, -0.0426326, 0.0746986, 0.1261370, 0.0710417, -0.1131095, 0.1187804, 0.1777732, -0.0826669, 0.1004176, -0.0594305, 0.1263376, 0.1975911, -0.1067853, -0.0571265, 0.1482562, -0.0251760, 0.1548684, -0.0057110, 0.0849441, 0.0044595, 0.1928194, 0.0745662, -0.0749171, -0.1340008, 0.2033060, -0.1515315, 0.1951771, 0.1295950, 0.0363555, 0.1166200, -0.1327413, 0.0487461, 0.0277203, 0.2546499, -0.1542276, -0.0682421, -0.1338578, 0.0697413, 0.4252724, -0.0396298, 0.0826924, -0.4392492, -0.2062666, -0.0481004, 0.3060647, 0.1037591, -0.0375688, 0.3107632, -0.1468026, -0.5094826, 0.2200745, -0.2497051, 0.2991661, -0.0216667, -0.0917714, 0.6292161, -0.0591128, -0.0071552, 0.1175462, -0.3466365, -0.4298849, 0.1137112, 0.2412775, 0.1082352, 0.0192067, 0.1291292, -0.1906887, 0.1214044, 0.4111048, -0.0323212, 0.0024477, 0.0046326, -0.2104903, 0.2206837, 0.2743008, -0.2028640, -0.0044374, -0.0640850, 0.5507017, 0.2758949, 0.1298936, -0.1320965, 0.0149061, -0.0805456, -0.1372381, 0.3141145, 0.3078074, -0.0114149, -0.3330400, -0.3103126, 0.1344222, 0.1206267, -0.0215327, 0.0146178, 0.3541521, -0.0069324, -0.1880898, 0.0842152, 0.4217070, -0.3227427, -0.2847326, 0.2162779, -0.0035071, -0.2422750, -0.0713898, -0.1295616, 0.2553110, 0.0320803, -0.1213197, -0.0083882, -0.0339394, 0.0177707, 0.0044480, -0.0010368, -0.0096005, 0.0288189, -0.0322330, 0.0035982, -0.1354144, -0.0982022, -0.0157425, 0.0033070, 0.0159032, 0.0222779, 0.0034406, -0.0947038, -0.0271617, -0.0288706, 0.0408339, -0.0185667, -0.0889987, -0.0072446, -0.0056528, -0.0091551, -0.1327057, -0.0338491, 0.0076566, 0.0072557, -0.0237218, 0.0069854, -0.0236838, -0.0856615, 0.0015117, -0.0149409, -0.0521846, -0.0064793, -0.0284085, 0.0867202, -0.0476118, -0.0094237, -0.1461497, 0.0281875, 0.0989131, 0.1315703, 0.2364842, -0.0523612, 0.2032122, 0.0131110, -0.0085451, 0.0780434, 0.0259757, 0.0735025, 0.0162738, -0.0627540, 0.0354236, -0.1070506, 0.1550144, 0.2168104, 0.1353535, -0.0008210, -0.0666923, -0.0590120, 0.0930269, 0.1937134, 0.0470727, 0.0805188, 0.1871244, 0.1566373, 0.0773064, 0.1948298, -0.0874235, -0.0354339, 0.1068951, -0.1227802, -0.1463703, 0.0749884, -0.0058918, -0.0469191, 0.3577731, 0.0821682, 0.0765989, -0.3383988, 0.1075600, 0.0512537, 0.0563210, -0.3823692, -0.0456547, 0.2011093, 0.2493168, 0.1375887, 0.0513697, -0.0143399, 0.0765535, 0.0038405, -0.0791382, 0.2901671, 0.0710372, 0.0234331, -0.2367113, -0.3706972, 0.1202276, 0.1072487, 0.0187939, -0.0392165, 0.1829972, 0.1497694, -0.0119939, -0.0278707, 0.2171601, -0.2475945, -0.0283204, 0.0620849, 0.0365405, 0.1258827, 0.1347727, 0.0326726, 0.0946533, 0.1082262, 0.2289364, -0.0285263, 0.0495861, -0.3018468, -0.1131763, 0.1709175, 0.1624923, -0.1989131, -0.0217438, 0.1881720, 0.0515522, 0.2065311, 0.0584583, 0.0979458, 0.1513012, -0.0129026, 0.1266432, 0.1005653, 0.0419965, -0.0673682, -0.1579996, -0.3605672, 0.1033390, 0.1347905, 0.1256807, 0.0363974, 0.2196113, 0.1689212, -0.0101414, -0.0428931, -0.0141052, -0.2033056, -0.0075726, -0.0539951, 0.0053848, -0.1147570, 0.1124537, -0.0193292, -0.0267614, -0.0405360, 0.1598528, 0.0285530, 0.1283026, -0.2063748, 0.0424266, 0.0458618, 0.0736743, -0.1661808, -0.0597049, 0.0215949, 0.3851948, 0.0930790, -0.0142903, -0.1239882, 0.0006748, -0.0434047, -0.1199295, 0.1314377, -0.0071033, 0.0238339, -0.2904101, -0.2836272, 0.1669919, 0.0344136, 0.0699019, -0.0686393, 0.0802572, 0.1537376, 0.0424847, -0.0009102, 0.2221003, -0.2921791, -0.0168269, 0.0734580, 0.0184599, 0.0499660, 0.1490703, 0.0467941, 0.1318561, 0.0216168, -0.2893601, -0.0341282, 0.0111168, 0.0060174, 0.0445205, -0.0257537, 0.0048543, 0.0603788, 0.0066666, 0.0191376, -0.1397964, -0.0532300, 0.0206533, 0.0328044, 0.0340700, 0.0275656, 0.0733631, -0.3200173, -0.0462968, 0.0253461, 0.0000928, 0.0288949, -0.0778521, -0.0028602, 0.0440229, 0.0093627, -0.2144318, -0.0094395, 0.0279379, 0.0160242, -0.0327548, 0.0200444, -0.0045957, -0.0917047, -0.0580307, 0.0107626, 0.0016237, -0.0071826, -0.0751732, 0.1056846, -0.1760277, 0.0800190, 0.0321362, 0.0734446, 0.0029748, 0.1188572, 0.1056639, 0.0814528, 0.0487020, 0.0094015, 0.0134020, -0.0675671, 0.0333399, 0.0423414, 0.0116104, 0.0337779, 0.1388162, -0.2755540, 0.0517918, 0.1833632, 0.0965308, 0.0159025, 0.0426725, -0.2719468, 0.1443281, 0.1541794, -0.1780030, 0.1894604, 0.0183333, 0.0562063, 0.0383339, 0.0897422, -0.0767570, 0.0503060, 0.1296381, 0.1434746, 0.0103961, 0.0401869, -0.0506201, 0.0651943, 0.3265342, 0.0585087, -0.0473572, -0.1824152, -0.2180606, 0.1968881, 0.1956099, -0.2244541, -0.0205022, 0.0071632, 0.2405656, 0.3060237, -0.0181665, -0.0904498, 0.1320747, 0.0660992, -0.0885849, 0.1790951, 0.2857963, -0.0684233, -0.1200168, -0.3243183, 0.0334017, 0.1422143, -0.0639363, 0.0493061, 0.2955657, -0.0028910, -0.0906863, 0.1158622, 0.1154760, -0.1380458, -0.1075904, -0.0162973, 0.0565629, -0.2857176, 0.0228605, -0.0116213, 0.1473116, 0.0872804, -0.0531366, 0.0341535, -0.1973920, 0.0119409, 0.0702701, 0.1582194, 0.2854652, 0.0570899, -0.0028334, 0.0457052, 0.3083474, 0.0794983, 0.1486394, 0.0241930, -0.2334183, -0.0749118, 0.2629755, -0.1049160, -0.0622753, 0.1039692, -0.1507371, -0.1539039, 0.0594115, -0.2021681, 0.2667516, -0.0349592, -0.0435668, 0.3692922, -0.0701067, 0.0074866, 0.2043889, -0.0345353, -0.3767520, -0.0315044, 0.0216058, 0.1653667, -0.1428512, 0.1308033, 0.0103670, 0.0089215, 0.2809844, 0.1460035, -0.0414160, 0.0490915, 0.0625192, -0.0083561, 0.0767171, 0.0578391, -0.0456690, 0.2480382, 0.2480070, 0.0509690, 0.0940972, 0.0555320, 0.0923206, 0.1828826, -0.1720205, 0.2568383, 0.1407311, 0.1187446, 0.0632933, -0.0309599, -0.0911574, 0.0128291, 0.0882619, -0.0106757, 0.2086174, 0.0499672, -0.0929909, 0.0865959, 0.2182694, -0.0396979, -0.0152263, 0.0010586, 0.0594860, -0.0337221, -0.0327425, 0.0552915, 0.0829210, 0.0010597, -0.0396099, 0.0282747, 0.0255513, 0.0029419, 0.0231883, -0.0762699, -0.0269072, 0.0212315, -0.0515209, -0.0084044, -0.1346324, -0.1271722, -0.1049417, -0.0138035, 0.0048985, 0.0337437, -0.0311930, -0.0474373, -0.0262088, -0.0500037, -0.0025950, -0.0377071, -0.0778910, -0.0727503, -0.0223368, -0.0810914, -0.1701600, -0.0529790, -0.0143296, 0.0100226, 0.0083356, -0.0146991, -0.0118568, -0.0671305, -0.0401891, 0.0061594, 0.0126762, 0.0176102, -0.0029477, -0.2474706, -0.0298180, 0.0815526, 0.1158801, -0.1637810, 0.0287815, 0.1376508, -0.0424984, 0.0670355, 0.2234169, 0.0213152, -0.0358289, 0.0337486, -0.0718430, -0.1614425, 0.0090935, 0.0828730, 0.0084185, -0.0881557, 0.2136187, 0.0087969, 0.1777235, 0.0439929, 0.0391467, 0.1755710, -0.0838418, 0.1634140, -0.0374354, -0.0267973, 0.1643859, 0.0187899, -0.1503244, 0.1672165, 0.1528651, -0.0518075, 0.0206415, -0.1065830, 0.1310139, -0.0916939, 0.1405271, -0.2316685, 0.2426717, 0.0633098, 0.1209891, -0.4417193, 0.1683812, -0.0069941, 0.0086475, -0.4441966, -0.0611136, 0.1705404, 0.4862059, 0.1423794, -0.0184582, -0.1627430, 0.0440884, 0.0010987, -0.2551653, 0.4215420, 0.0903071, 0.0509132, -0.1555232, -0.3586398, 0.1168805, 0.1141560, -0.0624483, -0.0366811, 0.1241965, 0.2147216, 0.0616217, -0.0188561, 0.3843378, -0.1690107, 0.0449388, 0.1051046, 0.0470401, 0.0465893, 0.1861739, -0.0146437, 0.1268283, 0.0628690, 0.1883257, 0.0695484, 0.1459658, -0.0491053, 0.0086274, 0.0730306, 0.1461562, -0.0045777, 0.0233239, 0.0175654, 0.0520265, 0.1229947, -0.0118564, -0.0066915, -0.0287755, -0.0340634, 0.2333643, 0.1138980, 0.0586095, -0.0417824, -0.1713802, -0.1798949, 0.1047944, 0.0382624, 0.0953299, -0.0060921, 0.0852891, 0.1361020, -0.0560700, -0.1069122, 0.1467122, -0.1030060, -0.0352063, 0.0857617, 0.0863729, 0.0946139, 0.1309477, 0.0329418, 0.1777034, 0.0614511, -0.0035876, -0.0427274, 0.0275480, -0.0403442, -0.0873260, 0.1329480, 0.1236226, 0.0247482, -0.0351283, 0.0413382, 0.3010016, 0.1248928, 0.1204591, -0.0687152, -0.0239718, -0.0490698, 0.0768626, 0.0946058, -0.0470454, 0.1183995, 0.0640410, -0.0435111, 0.1308724, 0.1230941, 0.2137360, 0.0951545, 0.0537363, 0.1947454, 0.0683797, -0.0695136, 0.0887816, 0.0023514, 0.0634278, 0.0975575, 0.1106803, -0.0369075, -0.0596941, -0.0153948, 0.0368063, 0.0005799, -0.1364068, -0.0729860, 0.0260791, -0.0081773, 0.0574077, -0.0262015, -0.0216833, 0.0653556, 0.0265399, 0.0030499, -0.1408897, 0.0202249, -0.0191565, 0.0567976, 0.0419143, 0.0322628, 0.0709652, -0.1788381, -0.0394902, -0.0331430, 0.0420086, 0.0798316, -0.0863712, 0.1185316, -0.0181413, -0.0112676, -0.1805472, -0.0459993, 0.0107849, -0.0251449, -0.0596815, 0.0629651, 0.0721377, -0.1144785, -0.0721719, -0.0129910, 0.0383648, -0.0346268, 0.0189326, -0.0438132, -0.0740595, 0.1377119, 0.2987877, -0.0818753, -0.0986169, 0.1918462, 0.0712813, 0.1394955, 0.2073626, -0.0068293, -0.1891705, 0.1640775, -0.1146807, -0.0302659, 0.0787281, 0.0541346, 0.2212257, -0.2669898, 0.1318246, -0.1932022, 0.2355520, 0.1529321, 0.0328492, 0.1405576, 0.0391682, 0.2864557, -0.0010477, -0.0817598, 0.0995812, -0.0787570, -0.1210288, 0.2183150, 0.1354482, -0.0488237, 0.1484968, -0.1302814, 0.1725622, -0.0465313, 0.2005635, 0.1083660, 0.1897793, 0.0696192, -0.1659742, 0.0077389, 0.1217660, 0.0060305, 0.1704886, 0.0973087, 0.0109273, -0.1020312, 0.2579273, 0.0533168, -0.0901949, 0.1037634, -0.0335824, 0.0488990, 0.0940165, 0.2077934, -0.0284255, 0.0246202, -0.1809940, 0.1226532, -0.0952619, -0.2528053, 0.0539649, -0.1052419, 0.2228697, 0.0995708, -0.2707940, 0.0399238, 0.2320437, -0.0492022, -0.1944864, 0.0598768, -0.0582705, 0.1810232, -0.1621256, 0.1589994, 0.1999080, -0.0115642, -0.0194252, 0.0738454, 0.0355164, -0.0292950, 0.1048165, 0.1479424, 0.2649528, 0.1546886, 0.2156552, 0.0058254, 0.1799057, 0.1166127, -0.0323718, 0.0478464, -0.0932458, 0.0050648, 0.3599487, -0.1567109, -0.0019182, -0.0194083, 0.0242839, 0.1134932, 0.0161761, -0.0111788, 0.1325444, 0.0061178, -0.0618391, 0.1444948, -0.0050981, -0.0531779, 0.1545531, 0.1504598, -0.0087875, -0.0808374, 0.1002335, 0.0775467, -0.0028395, 0.2352402, 0.1600343, 0.1800912, -0.1153438, 0.0221751, -0.1300231, 0.2363796, 0.1110382, -0.0439855, 0.0263370, 0.1563060, 0.1618621, 0.0093197, 0.2022138, -0.1612949, 0.1295603, 0.1639862, 0.0407651, 0.0968837, 0.0033178, -0.0292471, 0.1235911, 0.2318707, 0.0984067, 0.2020389, -0.0448425, -0.0460749, 0.0227461, 0.1035328, -0.1026051, -0.0076027, 0.0483123, 0.1281984, 0.0984853, 0.1409166, 0.0617327, 0.0744913, 0.0670084, 0.0924017, -0.1564923, 0.0566870, -0.0362449, -0.0468338, -0.2352235, 0.0216607, 0.0685882, -0.0859816, -0.0247470, -0.0744708, -0.0461078, 0.0281191, -0.0337683, -0.0984560, -0.2251123, -0.0635959, -0.1532766, 0.0061733, -0.0883845, -0.0289952, 0.0671707, -0.1657148, -0.0274146, -0.1449332, -0.0261116, 0.0461348, -0.0447968, -0.0437021, -0.0080223, -0.1202454, -0.2564536, -0.0968761, -0.0380930, -0.1120101, -0.1430482, 0.0265487, 0.0713491, -0.0587854, -0.0324532, 0.0212014, 0.1007260, -0.0309284, 0.0213873, -0.4062501, 0.0305455, -0.2316791, -0.0131648, -0.2795975, 0.1478137, 0.0091868, -0.1155339, 0.1177440, 0.2007220, -0.0506139, 0.1167569, 0.0933067, 0.1633348, -0.1668030, -0.1506414, -0.1527115, -0.0068280, 0.1960281, 0.0840781, -0.0977233, -0.0129105, 0.1761447, 0.2302029, 0.3031171, -0.2900133, 0.0298595, 0.0206465, 0.0211371, -0.2716255, -0.2529015, 0.1074125, 0.1919676, 0.0573884, 0.4383489, -0.2596429, 0.2620859, 0.1074997, -0.1294236, 0.1575466, -0.3868718, 0.1997886, 0.1061733, -0.0146264, -0.2264272, 0.2466503, -0.2008684, 0.0978202, -0.1953207, -0.1403699, 0.1975263, 0.4491968, 0.0297570, 0.1117057, -0.1169162, 0.0769187, 0.0236948, -0.2899092, 0.4830691, 0.1421883, 0.1060950, -0.1727753, -0.1280289, 0.0668442, -0.0483917, -0.1731638, -0.2906344, 0.2466133, 0.1572727, -0.0522876, 0.0013271, 0.3389462, -0.0617114, -0.0153503, 0.1182784, 0.0331060, 0.1204620, 0.0772107, 0.0693873, -0.0254149, 0.0776623, 0.1075735, 0.0962659, 0.0807748, -0.0712338, 0.1487759, 0.1063986, 0.0831166, 0.0104612, 0.0397779, 0.0709638, 0.2874934, -0.0061698, 0.0262751, -0.0179908, -0.0777962, -0.0539695, 0.1293582, 0.1789896, 0.1186673, 0.1159568, -0.0833234, 0.0015248, 0.1525858, 0.0663566, 0.1752154, 0.0053924, 0.1504938, 0.2465575, 0.0582539, -0.0728321, 0.3088160, -0.0165583, 0.0239112, 0.0469083, 0.1559511, 0.0776390, 0.0562722, 0.0861264, 0.1338668, 0.0960402, 0.0500441, 0.1936446, -0.0334219, 0.0080587, 0.1252470, 0.0097052, 0.0221647, 0.0955102, 0.0197011, -0.0298245, 0.1151668, -0.0373982, -0.1838017, -0.1018631, -0.0364622, 0.0342790, 0.1501189, 0.0659543, 0.1569855, 0.2585381, 0.1204419, 0.0842058, 0.0784548, -0.2082167, 0.0343740, 0.0524229, -0.1105358, 0.1498532, -0.0693922, 0.0681855, 0.2429806, 0.0426955, -0.1267756, 0.0236523, 0.4538180, 0.0283528, 0.0383992, 0.2568578, 0.1999253, -0.1597676, 0.0078541, 0.0132523, 0.2601731, -0.2072301, 0.0910817, -0.0169792, -0.1705959, -0.1434928, -0.1665801, 0.0687329, -0.1844618, -0.0966114, -0.2756105, -0.1316712, 0.0077918, -0.0955818, -0.0654567, 0.0810496, -0.0512312, -0.1515892, 0.0375422, -0.0181002, 0.1488179, 0.1831082, -0.0377191, -0.1550583, -0.1727127, 0.0023319, 0.0651674, -0.0904822, -0.0349028, 0.0621457, 0.1223454, -0.0207093, 0.0687098, 0.0035135, 0.2593353, -0.0884432, 0.1138168, -0.4275845, 0.0129906, -0.0423243, 0.3900101, -0.4690924, 0.1335146, 0.2043107, -0.0689861, -0.1740803, 0.1107772, 0.1702041, -0.1541852, 0.0948904, -0.2959923, -0.1411335, 0.0858735, -0.1190904, 0.2599701, 0.0408556, 0.1366097, -0.3226345, 0.1383294, 0.1810208, 0.3721279, 0.2064458, -0.1014637, 0.0061287, -0.0361531, 0.0574619, 0.0942447, -0.1552954, -0.0803286, 0.3031432, 0.2394475, 0.1935945, 0.3507061, -0.0594696, 0.4003660, -0.0963401, 0.1587182, 0.1177339, 0.0330266, 0.0634282, -0.0656258, 0.1139640, 0.0146071, -0.0116426, 0.0666491, 0.0984979, 0.1187969, -0.2520188, 0.1927238, -0.1100779, 0.1086255, 0.0533999, -0.0847456, 0.0275649, 0.1673165, 0.1599403, -0.0070922, 0.0369340, -0.2311994, 0.0903533, -0.0077260, -0.2708882, 0.0661687, -0.0264020, 0.1018603, -0.0627185, -0.1605354, 0.1144191, 0.0863379, -0.0274319, -0.0691343, 0.1795797, -0.0689749, 0.2095006, -0.0022345, 0.1431508, 0.1038172, -0.2130968, -0.1456293, 0.0022726, 0.5564734, -0.3641019, -0.0923098, 0.2858027, 0.0148664, -0.1509497, -0.1486277, 0.1968568, -0.1782844, 0.1924456, -0.3016339, -0.2943732, -0.0138525, -0.1740499, 0.5795859, -0.2111115, -0.0863535, -0.2537323, 0.0938611, 0.0236541, 0.5172631, 0.4140640, 0.2250903, -0.1416729, -0.2148384, 0.1760243, 0.3536924, -0.1559333, -0.1835051, 0.0979354, 0.2421430, -0.0799280, 0.3098370, -0.3120431, 0.6167250, -0.1778834, 0.0676789, 0.1634050, -0.2087064, -0.0440885, -0.0436244, 0.1780408, -0.0380081, 0.0294880, 0.1059029, 0.0938760, 0.1336087, -0.0267176, 0.0215360, -0.0216465, 0.1414872, 0.1443982, 0.0403239, 0.0282530, 0.0226646, -0.2328619, -0.0019109, 0.0817417, 0.0465027, 0.0816334, -0.0166346, -0.0620436, 0.0566603, 0.0988346, -0.1414514, -0.0132508, 0.1257847, 0.0864409, -0.0237283, 0.0250527, 0.0744061, 0.0217155, -0.0224590, 0.0286494, -0.0495561, 0.0375983, -0.0552733, -0.1741049, -0.1000395, -0.0539281, 0.2414826, -0.1546779, -0.0115227, 0.0332847, -0.2111191, -0.0444135, -0.0376163, -0.1592947, -0.1287573, -0.0327253, -0.1457217, -0.1393196, -0.3772884, -0.1135741, 0.0914184, 0.0620370, 0.0033994, -0.2961251, 0.0039374, 0.1125079, 0.2804636, 0.3225473, -0.0996886, -0.1162643, -0.0548270, -0.0984506, 0.0129519, -0.3160180, -0.0784357, 0.0781998, 0.2321972, 0.1529804, 0.0106319, 0.0442672, 0.2992834, -0.1586557, 0.1588139, -0.1907222, 0.1259561, 0.0118268, 0.0786720, -0.2652222, 0.1332663, -0.0744763, -0.0334800, 0.0256500, 0.0153951, 0.0030769, -0.0690117, 0.1181275, -0.1775932, 0.0236145, -0.1914690, -0.0518296, 0.0835694, 0.0462274, 0.0031001, -0.1283650, 0.0622292, 0.2080562, 0.1902105, 0.3527352, -0.3317888, -0.0925755, 0.0470367, -0.0543285, -0.0827896, -0.1267951, 0.0965078, 0.1889189, 0.0528000, 0.3410636, 0.0382944, 0.1039080, 0.1423700, 0.0662003, 0.1911118, -0.0901856, 0.2832746, 0.0033217, -0.1046117, -0.1347674, 0.0591361, 0.0107005, 0.1531257, 0.0404504, 0.0107610, -0.1528309, 0.0078340, 0.0349806, 0.0191207, 0.0842896, -0.2359970, -0.0864058, 0.0142803, 0.2410074, -0.1875199, -0.1927990, -0.2428914, 0.0469132, 0.1165348, 0.0553409, -0.2009584, -0.1153005, 0.1187260, -0.0697165, -0.3043111, -0.1640735, 0.3565593, -0.1660307, -0.2161292, 0.3077581, -0.1604229, 0.3828252, 0.0095799, 0.2314805, 0.2471315, 0.1381531, 0.0251801, -0.0335590, -0.0771436, -0.0061128, 0.1183147, 0.0625994, 0.1026823, 0.0750464, 0.0632707, 0.1857560, 0.1193456, -0.1474018, 0.2625239, 0.1812860, 0.2487425, 0.1300333, 0.1325279, 0.0286893, 0.0515800, 0.2033409, 0.1227187, 0.0866455, -0.0455821, 0.0008942, 0.0329462, 0.0479159, -0.0795120, 0.1852184, 0.1384540, 0.0506147, 0.1592024, 0.1117931, 0.0552086, -0.0400833, 0.2055765, 0.0267071, -0.1005323, 0.0826937, 0.0184784, 0.2964435, 0.1520340, 0.1703015, -0.1400745, 0.1719576, 0.0380186, 0.1370423, 0.2252971, 0.0632972, 0.0908231, -0.0777151, 0.0486322, -0.0361588, 0.1112557, 0.1829800, -0.1168095, 0.0514933, 0.4030021, -0.1230373, -0.0735240, 0.1491240, -0.1660485, 0.0139417, 0.0886413, -0.3676294, 0.2044583, -0.0543117, -0.0355287, -0.0040007, -0.0485457, 0.0578437, 0.1422216, -0.0861676, -0.1662228, 0.0455584, 0.2702916, 0.0667749, 0.0334112, 0.2913922, 0.1494647, -0.1367658, 0.1632419, 0.0691435, 0.2201944, -0.1759857, 0.0457568, -0.0020513, -0.0589857, -0.1109446, -0.1119053, 0.1227445, -0.1471806, -0.2189113, -0.2096331, -0.0449131, -0.1070843, -0.0156370, 0.0409127, 0.1075554, 0.0105200, -0.0867376, 0.0135502, 0.0825260, 0.2026666, 0.1630382, -0.1896553, -0.0612313, 0.0435382, -0.0197347, 0.0299669, -0.2331889, 0.0466785, 0.0243547, 0.2080103, 0.1048928, 0.1571839, 0.0672698, 0.2671955, -0.1402619, 0.2010929, -0.2086964, 0.0875638, 0.1311988, 0.3015586, -0.3769705, 0.1786020, 0.0831680, -0.2240234, -0.1312762, -0.0469836, 0.0258980, -0.2035522, 0.0068135, -0.4002886, -0.0525138, -0.0059777, -0.0352766, 0.2008667, 0.0241539, 0.0841508, -0.1665666, 0.0498206, 0.1982102, 0.2704237, 0.2634258, -0.2336503, -0.0504649, -0.0033806, 0.0274176, 0.0588252, -0.0131262, 0.1670048, 0.2045599, 0.2370483, 0.3171621, 0.2159330, 0.1228532, 0.3123582, 0.0713444, 0.2423526, 0.0674714, 0.0347805, -0.0717023, 0.0671098, 0.0438159, 0.0036248, -0.1018699, 0.1406012, 0.0635148, 0.0605209, -0.0947726, -0.0859249, -0.0140508, -0.0600522, 0.1373408, -0.1266407, 0.0040018, 0.0896969, 0.0454395, -0.0813947, -0.0217168, -0.1065172, 0.1318422, 0.0265575, -0.1578879, 0.0381401, -0.0937783, -0.0153442, -0.0995981, 0.0299576, 0.0328431, 0.0072462, 0.0512845, 0.0159066, 0.1477831, -0.1587241, 0.1385161, 0.1057880, 0.1169941, 0.0523420, -0.2008049, -0.1560530, 0.0436442, 0.5920684, -0.2848071, 0.0028922, 0.2969472, -0.3779324, -0.2892581, 0.0193054, 0.0661299, -0.1196468, -0.1006029, -0.3061673, -0.3290929, -0.1708928, -0.0604441, 0.2690352, -0.0090817, 0.1106803, -0.2125017, 0.1573142, 0.3268299, 0.5437714, 0.4853058, 0.0194783, -0.0766586, -0.2859329, 0.1354861, 0.2777056, -0.2030648, 0.0457190, 0.2142529, 0.4290656, 0.1856279, 0.3920025, -0.1005400, 0.6116643, -0.1281834, 0.2605555, 0.1480570, -0.0639408, -0.0817379, 0.0639149, 0.0887721, 0.0267681, -0.0500647, 0.0611473, 0.1136736, 0.0861188, -0.0053992, -0.1562165, -0.0633176, 0.1138792, 0.2292288, 0.0471647, 0.0492597, 0.1187128, -0.1508986, 0.0149639, 0.2074370, 0.0573299, 0.1507180, -0.0778908, -0.1049752, 0.0685572, 0.0438520, -0.2839581, 0.0763537, 0.1173652, 0.1694842, -0.0250421, 0.1475003, 0.1070818, -0.0320140, -0.0425557, 0.0399922, 0.0633565, -0.0039576, -0.0101465, -0.3038720, 0.0061435, -0.0833097, 0.4518305, -0.3957161, -0.0696592, 0.1074983, -0.1487300, -0.1730698, -0.0150657, -0.0762147, -0.2539669, -0.0788983, -0.2967061, -0.2598251, -0.2580340, -0.1716149, 0.0503802, 0.0589695, 0.0689261, -0.3100345, 0.1123897, 0.1210276, 0.5789589, 0.4527428, -0.0960075, -0.0477646, -0.0875706, -0.0217220, 0.2402166, -0.3110835, 0.0422297, 0.1464128, 0.2861869, 0.2370775, 0.1886557, -0.1119589, 0.4502024, -0.3508527, 0.1873265, 0.0408550, 0.1537936, 0.0951731, -0.0703632, 0.1165650, 0.0300043, 0.2474690, 0.1076539, 0.0165607, -0.0115436, -0.0431336, 0.2124980, 0.1358654, -0.0343569, -0.1320490, -0.0356854, -0.0447966, 0.0484913, 0.1336815, 0.1358303, 0.0943148, -0.1380347, -0.2621219, 0.1441873, -0.1577773, 0.1637468, 0.1201547, 0.1189091, 0.1286940, -0.0925455, 0.0290911, 0.0579057, -0.2662147, -0.1856804, 0.2671116, 0.1740415, 0.0728956, 0.0308735, 0.1133368, 0.1901667, 0.0824776, -0.1696078, -0.0348960, 0.0450809, -0.0445518, -0.0481611, -0.0204444, 0.0876901, 0.0553126, 0.0354004, -0.0031475, 0.0118563, -0.0407888, 0.0430293, -0.0181335, -0.0637519, -0.0561911, 0.0297962, -0.0347891, -0.0130740, -0.0458309, 0.0966315, 0.0462850, 0.0996111, -0.1089841, -0.0160096, 0.1175546, -0.1573183, -0.1125870, -0.0409956, -0.1085141, -0.1040352, 0.0676645, -0.0619919, -0.0817565, 0.0401024, 0.0462836, -0.0031465, 0.0370988, 0.0547041, 0.0040057, 0.1683275, 0.1335257, -0.0396098, -0.0250875, 0.0767314, 0.1820379, 0.1857133, 0.0048964, 0.0247522, 0.1399949, 0.1033769, 0.1976722, 0.1246421, -0.0641449, 0.0636339, -0.0221704, 0.0644883, 0.0702876, 0.0835788, 0.0632190, 0.0732044, -0.1335708, 0.0718395, 0.1973962, -0.0216354, 0.0294567, 0.1418305, 0.1996332, 0.0918254, 0.1375080, 0.1492884, -0.1322394, 0.0208232, 0.2661977, 0.0264112, 0.0216524, 0.0209160, -0.0528302, 0.1689374, 0.0108587, 0.0412543, -0.1688954, 0.1313013, -0.0310093, 0.0942226, 0.1756855, 0.1818446, -0.0131976, 0.2604378, -0.0513063, -0.0892099, -0.0205345, -0.1172721, 0.1261758, -0.0156166, -0.0282212, 0.3081245, 0.0378914, 0.0746645, -0.0263275, 0.0286066, 0.1243954, 0.1553971, 0.0270993, 0.0931610, 0.1904479, 0.0582928, 0.0407266, 0.1438244, 0.0526339, -0.0630046, 0.1433443, -0.0062140, 0.0999287, 0.0675981, 0.0069900, 0.1590123, 0.1841581, 0.2519496, 0.2347528, 0.2789993, 0.1499870, -0.0474945, 0.1224593, 0.1168787, 0.2694648, 0.1930118, 0.0699841, 0.1348860, 0.0146066, 0.3363145, 0.2037336, 0.0292028, -0.0658400, -0.0780902, 0.0372138, 0.1343911, 0.2537500, 0.2631676, 0.2207780, -0.2247405, -0.1726687, 0.1677050, -0.0648953, 0.2586871, 0.1113662, 0.3018071, 0.1268517, -0.0262322, 0.1524723, 0.2618069, -0.3629011, -0.2449483, 0.1923321, 0.1009024, 0.0798153, -0.0127784, 0.2673520, 0.2510564, -0.0299119, 0.0719267, -0.0407773, 0.0786283, -0.0681840, 0.0844204, 0.0857369, 0.1576364, 0.0192237, 0.0176083, -0.1089510, -0.0878256, -0.0325276, -0.2597482, -0.0989458, -0.0072629, -0.1561591, 0.1670569, 0.0544007, 0.1760383, -0.0969168, 0.0587472, 0.0494323, 0.0695357, 0.0218900, -0.0589445, 0.0110233, 0.1214624, 0.0446263, 0.0860018, 0.0266628, 0.0951895, 0.1766518, -0.0475157, 0.0229976, 0.1108357, -0.0305162, 0.0972950, 0.0477233, 0.2039696, 0.0014178, 0.2682229, 0.0236576, -0.1646305, 0.0952235, 0.1223386, 0.0330976, 0.1126866, 0.1535802, 0.1336425, 0.1449798, 0.2405610, 0.2315041, 0.1579964, 0.1201658, 0.0328975, 0.0781099, -0.0327502, 0.1517247, 0.2551198, 0.0724003, -0.0328687, 0.0670704, 0.0363173, -0.0200026, -0.0118674, 0.0986993, 0.3197023, 0.0125378, 0.0018045, 0.0450946, 0.2557816, 0.0689211, -0.0721909, 0.1298842, 0.0409621, -0.0900516, -0.1015775, -0.0122642, 0.2016265, -0.0354065, -0.0192455, -0.0227220, -0.0510347, 0.0515113, 0.1294750, 0.0623751, 0.1286789, -0.0171873, -0.0494513, -0.1123328, 0.1253105, -0.0509273, -0.1098425, -0.1033669, -0.1811182, -0.0880067, 0.0901485, 0.0641723, 0.0946944, -0.0129362, -0.0811015, -0.0876565, -0.0082162, -0.1080431, 0.0794604, -0.0033833, -0.0194054, 0.1240464, 0.0441999, 0.0617359, 0.1551571, 0.0327457, -0.0859782, 0.0280752, 0.0571210, 0.0306230, -0.0182013, 0.1215727, 0.1307101, 0.0260062, 0.3603401, 0.1293576, -0.1675354, 0.0030728, 0.1202725, 0.2142726, 0.1069673, -0.1342399, -0.1363375, 0.0606090, 0.3320417, 0.0911919, 0.0212969, -0.2037586, 0.0148741, -0.0158273, -0.0860646, 0.2508171, 0.2731049, 0.0082597, -0.2167179, -0.1718809, 0.0400661, -0.1665184, 0.0685436, -0.0301585, 0.1918756, -0.0709282, -0.2432912, 0.0992252, 0.2979211, -0.2921829, -0.1966905, 0.2700018, 0.0936553, -0.0615207, -0.0043396, 0.1590867, 0.2015952, 0.1876316, 0.1391036, 0.0465951, -0.0599274, 0.1462124, 0.0181870, 0.1884082, 0.1077471, 0.0385682, 0.0466025, 0.0030467, 0.1302958, 0.1028903, 0.0315407, 0.0741484, 0.0325134, 0.0125295, 0.0618709, 0.1093677, 0.1786675, 0.0902123, -0.2057989, -0.0449499, 0.1311821, -0.0696331, 0.1642020, 0.0376293, 0.1531096, -0.0030566, -0.0597077, 0.1364779, -0.0186006, -0.0840433, -0.0874931, 0.1570322, 0.0409188, 0.0355250, -0.0248068, 0.1237207, 0.1333321, 0.1493086, 0.0718218, 0.1543091, 0.0891441, 0.0294906, -0.0569477, 0.2246306, 0.0133281, -0.1104244, -0.1272486, -0.0142730, 0.3254014, 0.0456926, -0.0363078, -0.4497087, -0.0586925, -0.0291748, 0.0373853, 0.0892863, 0.1145844, 0.0794961, -0.1321125, -0.3441940, 0.1794273, -0.1569188, 0.2421591, 0.0294723, 0.1627199, 0.3158809, -0.0508919, 0.0109455, 0.1486796, -0.3753704, -0.2363046, 0.1422736, 0.2808909, 0.1004895, 0.1760261, 0.1156294, -0.0034639, 0.0682850, 0.2949685, 0.0811030, 0.0398897, -0.0849980, 0.1077577, 0.0561862, 0.2044023, -0.0629760, -0.0449571, 0.1873843, 0.0871787, 0.1304621, -0.1842661, -0.0117765, 0.0436062, 0.0509744, 0.2165757, 0.1757781, -0.0314659, -0.1201803, -0.1593925, -0.1084462, 0.1610490, 0.2075996, -0.1982922, -0.0382048, 0.3411678, 0.0439764, -0.1538070, -0.0962167, 0.1119223, -0.1346490, -0.1187095, -0.0438592, -0.0314539, -0.0960432, 0.1172192, 0.0949131, 0.1068963, -0.1891303, 0.4246079, 0.3254913, 0.0799883, -0.1572946, 0.2833700, 0.1300438, 0.1718702, -0.1940769, -0.0325843, 0.1934831, 0.4500311, 0.1364456, -0.0927435, -0.2759068, 0.1847270, 0.1016871, -0.1721620, 0.4349525, 0.2082500, 0.0896296, -0.1585984, -0.1183347, 0.0686600, 0.1814383, -0.0249750, -0.0686405, 0.3740884, 0.2405209, -0.2201842, 0.1191847, 0.4285695, -0.2642462, -0.1298507, 0.1723919, 0.2850176, 0.0698067, 0.1567911, 0.3166834, 0.3753047, -0.0211026, -0.0114510, 0.0711551, 0.0345044, -0.0695192, 0.0239874, 0.0081489, 0.0106700, 0.0138825, -0.0335933, 0.0238141, -0.0646076, -0.0276691, -0.0555720, -0.0350667, -0.0142715, -0.0142742, 0.0109894, -0.0119079, 0.0258533, -0.0312924, 0.0156359, -0.0059595, -0.0011453, 0.0282537, 0.0055403, -0.0643180, 0.0067322, -0.0226687, 0.0004763, -0.0419999, 0.0169585, -0.0033593, -0.0233460, -0.0814509, 0.0149742, -0.0547773, -0.0174978, 0.0054330, 0.0396291, 0.1379396, 0.0042040, 0.0569367, -0.1565075, 0.2171064, 0.0953598, -0.0045927, 0.0500970, 0.0663084, 0.0607633, 0.0683283, 0.2020705, 0.0275559, 0.1037649, 0.0993885, 0.0286520, 0.0979926, 0.1371379, 0.0292175, 0.1498795, 0.3074419, -0.0274716, 0.0573378, 0.1091288, 0.0023266, 0.1721239, 0.0514220, 0.0251566, 0.1490523, 0.1082108, 0.1445758, 0.0279016, 0.0184862, 0.0666148, 0.0795440, 0.1089106, 0.0237955, -0.1248874, 0.1374535, -0.0559262, 0.0171406, -0.1175288, -0.0688167, 0.0392874, -0.0104908, -0.0574992, 0.1044844, 0.0077227, -0.0138131, 0.0224439, -0.0805130, -0.1023592, -0.1062518, -0.1631327, -0.0580317, -0.0103649, -0.0606283, 0.1311944, -0.1370545, 0.1098532, -0.0554311, 0.0683799, 0.0588933, 0.0602250, -0.0164686, 0.0585916, 0.0154139, -0.0539383, -0.0225685, 0.0990113, -0.0125372, -0.0111526, 0.0766453, -0.0397520, -0.1198226, 0.1345881, -0.0400845, 0.0956226, 0.1078617, 0.0356733, -0.1231400, 0.5355052, 0.1885089, 0.0470606, -0.1653852, 0.3112031, 0.1443068, 0.1596534, -0.3256435, 0.0058497, 0.1204244, 0.6392979, 0.2009177, 0.0825878, -0.1585991, 0.1107547, 0.1032391, -0.2714382, 0.5184678, 0.4511772, 0.0820054, -0.1274612, -0.1405776, 0.0529274, 0.1059817, -0.0957141, -0.0113035, 0.4646340, 0.0771344, -0.2822644, 0.1398118, 0.3770774, -0.1281236, -0.0698600, 0.1465276, 0.1160939, -0.0474414, 0.0628624, 0.1746953, 0.4220108, 0.0922002, -0.0950853, 0.1453221, -0.0079616, 0.0602606, -0.1465178, 0.0048589, -0.1171366, 0.0694504, -0.1562640, -0.1607924, 0.1080490, -0.4113617, -0.1613809, -0.1628995, -0.1489200, 0.0138633, 0.0480095, -0.0223217, 0.0521668, -0.0021124, 0.0358755, -0.0735658, -0.0742601, -0.2542415, 0.1683819, -0.0021990, -0.2131882, -0.0731193, -0.1482046, 0.0691240, 0.0778150, -0.0625187, -0.0844744, -0.0044356, 0.1183387, -0.0299830, 0.0272424, 0.1492350, -0.0022619, 0.0579503, 0.3151160, 0.2563281, -0.0187562, 0.0436393, 0.0840626, 0.3109300, 0.1284917, -0.1150906, -0.0246699, -0.0168207, 0.4933045, 0.1150539, -0.1247757, -0.2027697, 0.1081201, 0.0536036, -0.1012236, 0.3857854, 0.2987896, 0.0987988, -0.3700193, -0.3886504, 0.0530863, -0.0194355, 0.0601770, 0.0249491, 0.3993015, 0.0383397, -0.2438171, 0.2434488, 0.3930179, -0.2681498, -0.2686526, 0.1203390, 0.3110208, -0.1351065, -0.0674640, 0.2491807, 0.2399382, 0.0426718, 0.0159397, -0.0106812, -0.0247903, 0.0403557, 0.0258749, 0.0099123, 0.0088832, 0.0052875, 0.0464713, 0.0046532, 0.0844160, 0.0650996, 0.0102650, 0.0198097, 0.0009217, -0.0115405, 0.0180114, 0.0396634, 0.0690885, 0.0502247, -0.0384941, -0.0347568, 0.0372335, -0.0086484, 0.0513967, 0.0774115, 0.0707678, 0.0321621, 0.0391028, 0.0619967, -0.0599703, 0.0206317, -0.0082504, 0.0410451, 0.0361720, -0.0633254, -0.0563719, 0.0383629, -0.0369609, 0.0045098, -0.1697123, 0.0840292, 0.0535259, 0.0375246, -0.1094207, 0.1908445, -0.0640831, -0.0594874, -0.1076179, -0.0223822, 0.1370844, -0.0705857, -0.0923148, -0.1744263, -0.1525162, -0.0579307, 0.2131040, -0.2077634, -0.0103921, 0.0652010, 0.0153381, -0.0333372, 0.2056730, -0.2238957, 0.1764861, 0.0324293, -0.1497787, 0.1873618, 0.0321924, 0.0434761, 0.0098639, -0.0501727, -0.0860106, -0.0037658, 0.2767101, -0.0934603, 0.1070644, 0.1599282, -0.2002296, -0.0059748, 0.3790264, 0.1051022, 0.1439842, -0.3945685, 0.0658274, 0.1857219, 0.0842087, -0.3015032, -0.1602307, 0.1766931, 0.2910487, 0.2481712, -0.0052962, -0.0207899, 0.1098591, 0.0090225, -0.0131505, 0.3109168, 0.0797069, 0.0029822, -0.3499309, -0.3383823, 0.1626797, 0.1008070, 0.0662538, -0.0785890, 0.2465461, 0.2012512, -0.1000680, -0.0083248, 0.2289190, -0.3311907, -0.0255997, 0.1038974, 0.0042791, 0.0579147, 0.1579538, 0.0921483, 0.1618512, -0.2611219, 0.6068956, 0.2343474, 0.0072907, -0.1788029, 0.2754397, 0.1701864, 0.2547791, -0.3506566, -0.1812105, 0.0385822, 0.5590577, 0.2686051, 0.0709729, -0.3165005, -0.1194895, -0.0567503, -0.1989221, 0.7080072, 0.2637437, -0.0366318, -0.4536475, -0.3193572, 0.1230983, 0.0082170, -0.2085143, -0.0566893, 0.4414335, 0.1948873, -0.3391539, -0.0480643, 0.5493568, -0.4240646, -0.3307157, 0.2987931, 0.0611840, 0.0423458, -0.0022099, 0.2009294, 0.4018497, -0.0168615, 0.0722998, 0.0565833, 0.0578198, -0.0280669, -0.0068225, -0.0005178, 0.0000572, -0.0108941, -0.0468859, 0.0363719, 0.0845327, 0.0383664, 0.0103966, -0.0016094, 0.0377527, 0.0421029, -0.0780719, 0.0855783, 0.0526290, -0.0023066, -0.0364045, -0.0405265, 0.0517951, 0.0826539, 0.0157084, -0.0242179, 0.0811683, 0.0295390, -0.0205635, -0.0050758, -0.0008482, -0.0619560, 0.0376658, 0.0282303, 0.0198865, -0.0285320, 0.0600970, -0.0071358, 0.0514882, 0.1785150, -0.2504534, -0.0010274, -0.2166580, 0.2270463, 0.0319546, 0.0584149, -0.0259312, 0.1467101, 0.1733550, 0.1230147, 0.0854546, -0.0356524, 0.1963008, 0.2001282, 0.0391920, 0.0988104, 0.0696249, -0.1609900, 0.0632137, 0.3316289, 0.1372642, 0.1662972, 0.0308685, 0.1695068, 0.0646250, 0.2299303, -0.1032467, 0.0622445, 0.1070228, 0.1237489, -0.0711257, 0.1449546, 0.1218873, -0.0152879, 0.0515174, 0.0347665, -0.2610798, 0.0355910, -0.1612162, 0.0852969, -0.2103738, -0.0029054, 0.0228954, 0.0418014, -0.0025687, 0.0713175, 0.0487959, 0.0447223, 0.0753329, 0.0103607, -0.1412525, -0.0412319, 0.0262874, 0.0407763, -0.0009342, 0.0006591, 0.1690879, -0.2182043, 0.0215215, 0.0036211, 0.0644626, 0.0491085, 0.0124208, 0.0100912, 0.0691394, 0.0631220, -0.1359826, 0.0035330, 0.0332113, 0.0267374, -0.0095643, 0.0371138, 0.0030362, -0.0229089, 0.0465685, 0.0068248, -0.0024611, 0.0407137, -0.0213041, -0.1709219, 0.5314544, 0.1989157, 0.1003266, -0.3825761, 0.0183543, 0.0679443, 0.1856344, -0.4823342, -0.1936453, 0.0625375, 0.4174999, 0.2337001, -0.1902625, -0.1924438, 0.1580267, 0.0153031, -0.1523976, 0.3798762, 0.1619632, -0.0925926, -0.3605045, -0.3868404, 0.1103479, 0.0487474, -0.1730902, -0.1759627, 0.3962051, 0.1557568, -0.1567558, 0.0261973, 0.2631463, -0.3447343, -0.1228176, 0.0146762, 0.1450779, -0.1228768, 0.1166462, 0.0950060, 0.3462633, 0.2713552, -0.1815543, 0.2075537, 0.0818369, 0.1926007, -0.2316712, -0.0139045, -0.0802729, 0.2184483, -0.0458327, -0.1846697, -0.0926998, -0.1639895, -0.1061359, 0.0640399, -0.0590519, 0.2161831, 0.2247206, -0.1940641, 0.0715690, 0.0070101, 0.0326860, 0.0834466, -0.0927730, -0.4201861, 0.0126334, 0.0095439, -0.2046016, -0.0865910, -0.1966625, 0.1072612, -0.1213732, -0.0892018, 0.0038532, 0.0780724, 0.0837613, 0.0540891, 0.0847655, 0.1369028, -0.0743658, 0.1358689, 0.4719633, 0.1260938, 0.1024726, -0.2069359, 0.0322106, 0.1384696, 0.2481380, -0.3134089, -0.3322294, 0.3044851, 0.3233216, 0.2376999, 0.0222406, 0.0785551, 0.2026780, 0.0055463, 0.0453039, 0.2291087, 0.0213064, 0.0599771, -0.4397986, -0.4013881, 0.2487824, -0.0006563, 0.1832236, -0.2581193, 0.3589427, 0.3726108, 0.0002733, 0.0411070, 0.1406486, -0.4845511, -0.2123096, 0.0112682, 0.0000890, -0.0371939, 0.2078680, 0.0585039, 0.0834977, 0.0031523, -0.0933497, -0.0288776, -0.0905438, 0.0143530, -0.0140302, 0.0145391, -0.0050801, 0.0044460, 0.0474478, 0.0074391, 0.0459036, -0.0589668, 0.0254467, -0.0212032, -0.0075207, -0.0170788, -0.0137874, -0.0741144, -0.0369815, 0.0439388, 0.0137603, 0.0014629, -0.0164928, -0.0120916, 0.0478754, 0.0349683, -0.0235614, 0.0141469, 0.0051437, -0.0068191, 0.0064937, 0.0281353, -0.0217620, -0.0645040, 0.0229425, -0.0407987, -0.1725939, 0.0128019, -0.0495925, 0.0947538, -0.4178009, 0.0502746, 0.0385797, 0.0903378, -0.0993143, 0.0401897, -0.0030202, 0.0695916, 0.0246334, -0.1384673, -0.1271030, -0.2058740, -0.1164778, 0.0425544, -0.1385648, 0.0313305, 0.3755128, -0.3572099, -0.0346268, 0.0197994, 0.0740536, 0.2260990, -0.0361682, -0.2392109, 0.0845845, 0.0344090, -0.2993772, -0.0359452, -0.0195241, 0.0273927, -0.0972287, 0.0885480, -0.0100647, -0.0459543, 0.0546730, 0.0185701, 0.0570890, 0.0940081, 0.0119179, -0.0540706, 0.3659184, 0.1282776, 0.0856394, -0.3482178, 0.1137138, 0.0162217, 0.0293593, -0.3625402, -0.0519321, 0.1440544, 0.3376085, 0.1788035, 0.0591614, 0.0155733, 0.1274960, 0.0617009, -0.2286008, 0.3605622, 0.0671716, 0.0022187, -0.3021542, -0.3307347, 0.0771594, 0.1537159, -0.0626782, -0.0450943, 0.2180102, 0.0928740, -0.0281982, 0.0011492, 0.2695649, -0.3111356, -0.0040268, 0.0654196, -0.0279764, 0.0216400, 0.1156609, 0.0090740, 0.1267631, -0.3089703, 0.5178255, 0.3367148, -0.0132748, -0.2847394, 0.2735174, 0.1098433, 0.1308836, -0.3104376, -0.1371694, 0.0348851, 0.8310027, 0.2801426, 0.0288253, -0.3234674, 0.0582086, 0.2176924, -0.3423816, 0.6138118, 0.2835157, 0.0343955, -0.5255246, -0.3853560, 0.0122109, 0.0677300, -0.1857951, -0.0047190, 0.3216711, 0.1091856, -0.4522457, 0.0570299, 0.6991123, -0.3640231, -0.1743529, 0.2036373, 0.2184169, -0.0109656, 0.1077192, 0.2091782, 0.4832528, -0.0580124, 0.2480334, 0.0229831, 0.0670625, -0.0905863, 0.0170443, 0.0447554, 0.0087336, -0.2830826, -0.0765067, 0.0994487, 0.1735181, 0.0589144, 0.0807200, -0.0067179, 0.0616073, 0.0230395, -0.3349654, 0.2417058, 0.0278795, 0.0182129, -0.1079252, -0.2614173, 0.1213893, 0.0547276, -0.0487971, -0.0012385, 0.1468520, 0.0638360, 0.0832027, 0.0146014, 0.1230588, -0.2875471, 0.0494451, 0.0844639, 0.0354003, -0.0833711, 0.0619929, -0.0464862, -0.0002943, -0.0132816, 0.0214492, -0.0165319, -0.1458586, 0.1966829, -0.0522590, -0.0377473, -0.0890883, 0.1541976, 0.1216744, 0.0711655, 0.1153477, -0.0687564, 0.1704688, 0.2017749, 0.0553051, 0.0820424, -0.0512406, -0.0321558, 0.0476383, 0.1517569, 0.0387000, 0.1915935, -0.0486096, 0.0335382, -0.0330299, 0.0697194, -0.0114877, 0.0004333, 0.0010810, 0.0940928, -0.0711892, 0.1152685, 0.0904363, -0.0091679, -0.0351201, 0.0027588, -0.1446795, 0.0067526, -0.1259345, 0.0903798, -0.0430143, 0.0218382, 0.0444137, 0.0394465, 0.0112501, 0.0256840, 0.0846999, 0.0849275, 0.0324478, 0.0383828, -0.1012682, 0.0531193, 0.0233835, 0.0795208, 0.0098272, 0.0602253, 0.1063683, -0.1059586, 0.0137202, 0.0165438, 0.0488062, 0.0346676, 0.0460355, 0.0368570, 0.0271571, 0.0468416, -0.0493314, 0.0044588, 0.0338430, 0.0146836, 0.0174050, 0.0350957, 0.0415239, 0.0186603, 0.0152364, 0.0426590, 0.0370546, -0.0007953, 0.0070369, -0.0177405, 0.1685227, 0.0281002, -0.1530763, -0.0607477, 0.1192492, -0.0491943, 0.0990404, 0.0138339, -0.0379554, 0.1708068, 0.2986441, 0.0830394, 0.1196502, 0.0746222, 0.0937407, 0.0478573, -0.0587780, 0.2299557, 0.0072108, 0.1246672, -0.1558541, -0.1093395, -0.0453323, 0.0211310, 0.1176149, -0.0430805, 0.1388868, 0.0938648, -0.0531083, 0.0818820, 0.1064282, -0.0519832, -0.0689414, -0.0109739, -0.0395969, 0.0166844, -0.0724576, 0.0694818, 0.0105536, 0.1954732, -0.0218400, 0.2170451, 0.2410814, 0.2337825, -0.0738998, -0.0027692, 0.1193743, 0.2695830, 0.0492394, -0.1307545, -0.1314358, 0.0442262, -0.1865164, 0.4443254, -0.1096803, 0.1643705, 0.2139710, -0.1654271, 0.0655322, -0.1101799, -0.1016381, 0.2421872, 0.1166415, -0.2827991, -0.0913156, -0.0205920, -0.0320770, -0.1881713, -0.0556334, 0.0283199, -0.0308517, -0.0047393, 0.1751901, 0.2438177, 0.1414745, 0.2467112, 0.2937405, 0.0630096, -0.0796440, 0.0540497, 0.2746934, 0.1163357, -0.0426831, -0.0108241, 0.1317774, 0.0209482, 0.0078605, -0.0568676, -0.0245622, 0.2192285, 0.3178022, 0.1252632, 0.1742059, 0.0672436, 0.1547868, 0.1556024, -0.2479261, 0.2895662, 0.1502314, 0.1521203, -0.0708120, -0.2024857, 0.0137782, 0.2525128, 0.0781370, 0.0847931, 0.2045707, 0.1089979, 0.0480602, 0.0784250, 0.1554254, -0.1732475, 0.0717787, 0.0119614, -0.0361945, -0.0139201, -0.1021589, 0.0268240, -0.0387832, 0.0267436, -0.2090103, -0.0137610, -0.1127278, 0.0605683, -0.0218959, -0.0502859, 0.0006967, 0.0421813, 0.0141261, 0.0025351, 0.0018755, -0.1610675, 0.0092206, 0.0320481, -0.0015858, 0.0243700, 0.0132619, -0.1846748, -0.0295099, 0.0236013, 0.0370058, 0.0480332, -0.0870092, -0.0521453, -0.0074125, 0.0130600, -0.1784447, -0.0210977, 0.0225279, 0.0168592, -0.0186776, 0.0168626, -0.0052654, -0.0391723, -0.0091444, -0.0135828, -0.1537417, 0.0061022, -0.0652040, 0.1263169, -0.3643431, 0.0170790, -0.0019764, 0.0495796, -0.0647821, 0.0231456, -0.0111999, 0.0510630, 0.0489444, -0.1480415, -0.1869196, -0.1553259, -0.0503561, 0.1020452, -0.0078523, 0.0217372, 0.3401100, -0.3252890, -0.0040763, -0.0229599, 0.0151665, 0.1124922, -0.0593720, -0.2128415, 0.0481191, -0.0058960, -0.2723763, -0.0120674, -0.0282584, 0.0721126, -0.1034541, 0.0672930, -0.0338855, 0.0171952, -0.0815501, 0.0591684, 0.0328364, 0.0848740, 0.0225827, -0.0848798, 0.2246644, 0.0821767, 0.0353540, -0.2170315, 0.0900950, 0.0396275, -0.0303367, -0.3524975, -0.0823549, 0.1323073, 0.4989445, 0.0409824, 0.0703220, -0.1480542, 0.0224627, 0.0512453, -0.2606803, 0.3512332, 0.1329067, 0.0199689, -0.1123916, -0.3217358, 0.0885997, 0.0816272, -0.0552667, -0.0050162, 0.0875352, 0.1229674, 0.0441924, 0.0158962, 0.3165502, -0.1621452, 0.0218151, 0.1341836, 0.0337414, 0.0563569, 0.1421688, 0.0104334, 0.0333876, -0.1376542, 0.4323340, 0.2396287, 0.0607290, -0.0599313, 0.0220720, 0.1068949, 0.1107977, -0.0510220, 0.1219104, -0.0179161, 0.7416416, 0.1469480, 0.1350228, -0.1084552, 0.1534379, 0.2378175, -0.3109058, 0.5340213, 0.2603593, -0.0073719, -0.1993406, -0.1164143, -0.0391089, 0.0756348, -0.2151570, 0.0965009, 0.2934655, -0.0773626, -0.3033855, 0.0537706, 0.4921612, -0.2293288, -0.0562078, 0.1469331, 0.0859654, -0.0412326, 0.0145451, 0.0524719, 0.4046888, -0.2630724, 0.1409971, 0.0648238, 0.2255224, -0.3074340, 0.1028372, 0.0899597, -0.2115159, -0.5319832, -0.1072161, 0.2296880, 0.3387732, 0.1763027, 0.0270030, -0.4361921, 0.0309635, 0.0061911, -0.3083101, 0.2670833, 0.2335424, 0.0306433, 0.0560054, -0.2062085, 0.2449556, 0.1656870, -0.2769188, 0.0753938, 0.1553710, 0.1285151, 0.1991051, 0.0139611, 0.1978070, -0.0414585, 0.1743431, 0.2141029, 0.2126459, -0.0385448, 0.2699521, -0.0656116, -0.0176028, -0.0546311, 0.1240107, 0.1107264, -0.1857068, 0.1349868, 0.1029668, -0.0759438, -0.0342413, 0.0643768, 0.0942879, 0.0415695, 0.1524955, -0.0032176, 0.1422403, 0.1114412, 0.0344350, 0.1227296, -0.1589247, 0.1400556, 0.0885339, 0.1336691, 0.0468377, 0.1398502, -0.0560669, 0.0856719, -0.0778825, 0.0231485, 0.0485336, -0.0005165, -0.0695553, 0.0424885, 0.1107770, 0.1177571, 0.0236100, 0.0557647, 0.0145289, -0.0448823, -0.1452113, 0.0391446, 0.0047189, -0.0095054, -0.0681843, -0.0760902, 0.1043582, 0.0086060, 0.0947092, -0.0209333, 0.0095728, 0.0323286, 0.0071412, -0.0295927, -0.1833839, 0.0454857, -0.0729210, 0.0400834, 0.0081658, 0.0086889, 0.0492315, 0.0033266, 0.0239286, -0.0288851, 0.0574660, 0.0593996, 0.0537443, 0.0715772, 0.0184797, 0.0390316, -0.0931672, -0.0017859, 0.0652938, -0.0390517, -0.0007657, 0.0311596, 0.0860594, 0.0520700, -0.0340422, 0.0770791, 0.1421760, -0.0469462, 0.0170053, 0.0949611, -0.0566984, -0.0096147, -0.1538580, 0.1387391, 0.0790826, -0.0926924, -0.0047629, 0.0683548, 0.0474823, 0.0530087, 0.1226216, -0.0864260, 0.1478869, 0.1551975, -0.0007358, 0.0472642, -0.0639180, 0.0233376, 0.0182589, 0.1284930, -0.0062571, 0.0326662, -0.0117146, 0.0276850, 0.0464716, 0.0635186, -0.0449919, 0.0458106, 0.0237422, 0.0454131, 0.0287730, 0.0377682, 0.0260776, 0.0647337, -0.0145770, 0.1149632, -0.1378173, 0.0483268, -0.1226717, -0.0878852, 0.0374052, -0.0061958, 0.4144586, -0.1259560, -0.0281462, 0.1568162, 0.0003380, -0.0071307, 0.1925666, 0.0399400, -0.0630550, -0.1084500, -0.1899728, -0.0589324, -0.1626205, -0.0210974, 0.1238761, 0.0797283, 0.2989622, -0.2237088, 0.3006380, 0.1868754, 0.4086194, 0.3106743, -0.1319402, 0.2184908, 0.0306804, -0.0842817, 0.0498379, -0.1973841, 0.0649129, 0.2549534, 0.3584079, 0.3387897, 0.4368521, 0.0089726, 0.5013810, -0.1107408, 0.3654904, 0.0535149, 0.0473498, 0.0000162, 0.0577032, 0.0445216, 0.0901664, 0.0052091, -0.0444381, -0.0852024, 0.0460915, 0.2095148, 0.1789627, 0.0333307, 0.1871535, 0.1673292, 0.0452259, 0.1158809, -0.3035533, 0.1224966, 0.1292208, 0.1195014, 0.1092280, 0.0373892, 0.1304447, 0.2286706, -0.0912825, 0.1312756, -0.0066113, 0.0849881, 0.1958906, 0.0557834, 0.1271151, 0.0662476, 0.2498266, 0.1436521, -0.0218035, 0.0264646, 0.0933849, -0.0931496, -0.1333767, 0.0442372, -0.1127347, -0.0227397, -0.0438933, 0.0376333, -0.0302466, -0.0282023, -0.0353642, 0.0561348, -0.0047426, -0.0004306, -0.1101222, -0.0867805, -0.0034159, 0.0358539, 0.0352031, 0.0188612, 0.0335232, -0.0738962, -0.0198958, -0.0278589, -0.0050822, 0.0268029, -0.0933032, 0.0361590, -0.0093115, -0.0140102, -0.1134880, -0.0364822, 0.0135144, 0.0174895, -0.0283853, -0.0136600, 0.0183916, -0.0442308, -0.0267276, 0.0090837, -0.0825713, -0.0141399, -0.0678271, 0.0228220, -0.3193049, -0.0353375, 0.1577225, 0.0154357, -0.0339672, 0.0403727, -0.0522699, 0.0591919, -0.0253615, -0.1331523, -0.1240624, -0.1508881, -0.1211916, -0.0464265, -0.0647958, -0.0360599, 0.0771842, -0.1568356, -0.0621653, -0.0820415, -0.0271787, 0.0390423, 0.1776482, 0.0007671, 0.0212921, 0.0235829, -0.2922193, 0.0502734, 0.0748925, 0.0239889, -0.0579365, 0.0211289, 0.0277717, 0.0319913, 0.0065487, 0.0446833, 0.1633697, 0.0125431, 0.1139461, 0.0573046, -0.0409477, 0.1430728, 0.0992092, 0.0587481, 0.0747174, -0.0190435, -0.1172358, -0.1116352, -0.0931931, 0.0292161, 0.2053453, -0.0965337, -0.0204631, -0.0616717, -0.0505910, 0.0977463, -0.0207149, 0.1160064, 0.0928131, 0.1318064, -0.0331050, -0.1017194, 0.0225174, -0.1191157, 0.0299139, -0.0349250, -0.0812816, 0.1253352, 0.0734560, 0.1744612, 0.0853463, -0.0894314, 0.0150194, 0.0455749, 0.1555886, -0.0889618, 0.0855090, 0.1399790, -0.1589440, 0.1245100, 0.3903219, 0.3917106, 0.0505790, 0.0618480, 0.1299539, 0.0639763, 0.0917409, -0.0771636, -0.0195120, 0.1797161, 0.5320565, 0.1100515, 0.0881272, 0.0775279, 0.3807711, 0.3781696, 0.0312439, 0.2743511, 0.2959478, 0.1664379, -0.0136636, -0.1599640, 0.0474853, -0.0709945, 0.0974605, 0.0017734, 0.4412239, 0.0216220, -0.0598408, 0.3440855, 0.3467680, -0.1009982, 0.0276164, -0.0452919, 0.2974166, -0.0823894, -0.0256282, 0.2747280, 0.1936014, -0.1202984, -0.0643450, 0.0907721, 0.1004114, -0.0165656, 0.2088750, 0.0659987, -0.0518615, -0.0484500, 0.0286073, 0.2920682, 0.0453509, -0.0557321, 0.0877433, 0.0290023, 0.0712988, 0.2169936, -0.1010760, 0.0436894, 0.2459426, 0.1276845, 0.1979513, 0.1157165, 0.2107936, 0.1936861, -0.1283235, 0.1747888, -0.0691280, 0.1091534, 0.1974754, 0.0006188, 0.1645447, 0.2264639, 0.3137963, 0.0615412, 0.3494515, 0.0397039, 0.2393015, 0.0078344, 0.0291937, 0.0560398, 0.1613093, 0.1966991, 0.0154676, 0.0307184, 0.1386042, -0.0307608, -0.0752767, -0.0305206, -0.0806119, 0.1287910, 0.1864278, -0.0407622, 0.0693999, 0.1358804, 0.1815882, 0.1831258, 0.0084790, 0.2573869, 0.1427400, 0.2078599, -0.0163818, 0.0358639, 0.0190881, -0.0226875, -0.0791543, -0.0323662, 0.0287056, 0.1049175, -0.0106627, 0.1141179, 0.1669583, -0.1190700, -0.0467716, 0.0748309, 0.2078396, 0.0598360, -0.0073629, 0.2133146, 0.0405413, 0.0100710, -0.1306457, -0.0167723, 0.2688087, -0.0698460, 0.0601051, 0.0749398, -0.1268988, -0.0299108, -0.0527685, -0.0735210, -0.1077266, -0.0262688, -0.2000283, -0.0221136, 0.0528011, -0.0055041, 0.0753912, -0.0777146, 0.1150815, -0.0681308, 0.1219836, 0.1102160, 0.1486188, 0.1537700, -0.0429787, -0.0494550, -0.2203990, 0.0184117, 0.1716735, -0.0517148, -0.0584696, 0.0301170, 0.1242514, 0.0327164, 0.1610131, 0.0016540, 0.1678636, -0.0075516, -0.0144158, 0.0668396, -0.2596839, -0.0346789, -0.0505285, 0.1055961, 0.0338849, -0.0310045, -0.0297662, 0.0386940, 0.0462688, 0.0122928, -0.0259500, -0.1096970, 0.1001358, 0.0874634, 0.0011748, 0.0267068, -0.0275489, -0.1513384, -0.0148521, 0.1214867, 0.0010852, -0.0129586, 0.0268082, -0.0520028, 0.0154760, 0.0497730, -0.2220086, 0.0745017, 0.0592119, 0.0343402, -0.0084529, -0.0249250, 0.0125192, 0.0441331, 0.0088006, 0.0500385, -0.0315710, 0.0372431, -0.1242334, -0.1774074, 0.2395493, 0.4032861, 0.1626290, -0.2629715, 0.3791557, 0.0902967, 0.0524597, -0.1503097, 0.0104695, 0.1656275, 0.2254258, -0.1145953, -0.2711464, -0.2832034, 0.1495066, 0.1106538, 0.2926292, 0.2692572, 0.5147160, 0.0691434, 0.0214942, 0.1214472, 0.2821761, -0.0261513, -0.1554965, 0.0507815, 0.1506738, 0.1368480, -0.0305626, -0.0098045, 0.3567445, 0.2250611, -0.0357590, 0.1540151, 0.6037115, -0.0098042, 0.2464386, 0.2638068, 0.4239621, -0.0138021, 0.0211125, -0.0076183, 0.2058673, 0.0647463, -0.0560189, -0.0223778, -0.0381489, -0.1420192, 0.0125520, 0.0440133, 0.0472521, 0.0114470, 0.1176926, 0.0972912, 0.1529854, 0.0156881, -0.0829540, 0.0200912, 0.1671085, 0.0185799, 0.0563110, 0.0262324, 0.1006765, 0.1626906, -0.0181751, 0.0774508, 0.0133418, 0.0777275, 0.2867609, 0.0859824, 0.0333271, 0.0280991, 0.2235091, 0.0977046, -0.0182532, 0.0064536, 0.1260903, -0.0585846, -0.0223196, -0.0700028, 0.0130481, -0.0301929, 0.1106490, -0.0402026, 0.0241549, -0.0355673, -0.1733747, -0.0587332, -0.0871696, 0.1103815, -0.1377438, -0.0351990, -0.1133109, 0.0140514, 0.0718044, -0.0191162, -0.0649991, 0.0748819, 0.0138008, -0.0900012, 0.0490287, 0.0616894, 0.0498753, 0.1189105, -0.0758488, -0.0536240, -0.0666714, -0.0361608, 0.0721163, -0.0483192, -0.0713020, 0.0688448, 0.0589384, -0.0782953, 0.0019855, -0.0399382, 0.0546158, -0.1085030, 0.0188585, -0.0462179, -0.0503578, 0.0026544, 0.2452643, -0.0824817, 0.1310730, 0.0629485, 0.0891295, 0.0745882, 0.1524707, -0.0996477, -0.1853585, -0.2364205, -0.1388036, -0.0322009, -0.0401999, -0.0059073, 0.1852531, -0.0601335, 0.0455726, -0.1108662, 0.1380788, 0.1773200, 0.2225219, 0.1117384, -0.0653084, 0.0745470, -0.2669076, 0.0293243, 0.2014904, 0.0263750, 0.0142781, 0.0782772, 0.2101665, -0.0184578, 0.0947117, -0.0159201, 0.3065294, -0.1282723, 0.0521751, 0.1612255, -0.2056130, -0.1508826, -0.0025471, 0.0930425, -0.1059792, 0.1656875, 0.1184453, 0.0608351, 0.0186264, -0.1450771, -0.0862469, -0.1477921, -0.0385804, 0.0139182, 0.0281424, 0.0319594, 0.1353673, -0.2187035, 0.0511988, 0.1035316, 0.0247788, 0.0416056, 0.1165266, -0.1015877, 0.1267367, 0.0761226, -0.1485055, 0.0379221, 0.2169207, 0.0625481, -0.1114222, 0.0496115, 0.1341871, -0.1078652, 0.0067754, -0.0137222, 0.1844191, 0.1172573, -0.0143939, 0.0300776, 0.0140790, 0.2616156, -0.0840939, 0.0654913, 0.1481141, -0.1062602, -0.0190207, 0.0528324, 0.0089270, 0.1643148, 0.0124191, -0.0576648, -0.0789676, -0.0175680, 0.0297905, 0.0309913, -0.1270936, 0.0547369, -0.0061077, 0.1047972, 0.0219670, 0.0554964, 0.0536887, -0.0926545, -0.0880381, -0.0059323, 0.0848406, 0.0719937, 0.0265839, 0.2103506, 0.0871884, 0.0498102, -0.0491656, 0.0255653, 0.2736609, 0.0477212, 0.0895085, 0.0708134, -0.0842386, 0.3081485, -0.1071337, -0.0319879, 0.0561971, 0.3659993, -0.1337974, 0.1145599, 0.0382633, 0.1997409, 0.2625251, 0.0104855, 0.0099589, -0.0420148, 0.3030824, 0.1783956, 0.1020506, 0.0110215, 0.0867876, -0.2049293, -0.0068352, 0.1104012, 0.1121377, 0.1236506, 0.1422863, 0.1130516, 0.0865090, 0.2161437, -0.1244666, 0.1208402, 0.2314815, 0.1303592, 0.0056523, 0.0706971, 0.1025841, -0.0464752, 0.0545848, 0.0667115, 0.0402444, 0.0500621, -0.0525851, 0.0338418, 0.1264974, 0.2744433, 0.0488093, 0.1729657, 0.0021172, -0.1027747, -0.0621526, -0.0288137, 0.0173664, 0.2576028, -0.0207553, -0.1230208, 0.1453763, 0.0365832, 0.2470388, 0.1856091, -0.0526991, 0.0761206, 0.0420395, 0.1471956, 0.1209147, 0.0713872, 0.0167037, -0.1146174, 0.0322944, -0.0256752, 0.0022067, -0.0239781, 0.0148948, 0.2958129, -0.0812481, 0.0008712, 0.1201529, -0.1706672, 0.1315265, -0.0768227, -0.0224999, 0.1383918, -0.0224630, -0.0278556, -0.0290996, -0.0147724, 0.2076365, -0.0028832, 0.0777688, 0.0496936, 0.0074878, 0.0441291, 0.1223077, -0.1008058, 0.0344444, 0.0186221, -0.0930835, 0.0498332, -0.0532454, 0.0816539, 0.2204410, -0.0264862, 0.1126825, -0.0015633, 0.1465884, 0.0868876, 0.0815501, 0.0623155, 0.0108345, 0.0535282, -0.0134929, -0.1400215, 0.1131136, 0.0505989, -0.0176536, 0.1071833, 0.0453197, -0.0815286, 0.1452297, 0.0168988, 0.2770569, 0.0500977, 0.1319232, 0.1190046, -0.0459477, -0.0667431, -0.0109100, 0.1908642, 0.0208246, -0.0200089, -0.0083040, 0.0391354, 0.0336377, -0.0078768, -0.0773990, -0.1707253, 0.1983444, 0.0603835, 0.0789586, 0.0617852, 0.0383397, -0.0246616, -0.0133348, 0.1584821, 0.0392746, 0.0013005, -0.0303015, -0.0261150, 0.0410652, 0.1624030, -0.2225479, 0.0422076, 0.1065500, 0.0928615, -0.0508319, -0.0075027, 0.0666495, -0.1252982, -0.0965287, -0.0360133, -0.0435690, -0.0633928, -0.0744363, -0.1093042, 0.1536993, 0.3495169, 0.0712008, -0.0473306, 0.3142379, -0.0537350, -0.0199192, -0.1815801, -0.1425466, 0.2870010, 0.1860696, 0.0153163, -0.2630615, -0.1243111, 0.0763169, 0.0606608, 0.1157200, 0.2858893, 0.2917948, 0.1375925, -0.0244130, 0.1565493, 0.0541894, 0.0574125, -0.1361913, -0.1783899, 0.0440546, 0.1087943, -0.0298720, 0.1549184, 0.2140271, 0.0705103, 0.1348353, 0.0436344, 0.3858768, 0.0857049, 0.2284125, 0.2410522, 0.2329329, -0.0945091, 0.2543360, 0.3098640, 0.1877653, 0.0142418, 0.2117128, 0.0095571, 0.0806612, -0.1453624, -0.0101585, 0.1257771, 0.1331818, -0.0989586, 0.0023420, 0.0057352, 0.0130669, 0.1965155, 0.1654590, 0.0583291, 0.2770292, 0.1740821, 0.1795466, 0.0417842, 0.0101734, -0.0013039, -0.0266102, -0.0339694, 0.0838667, 0.1105953, 0.1906180, 0.0056866, 0.2372436, 0.2061149, 0.1737709, 0.0118608, 0.3541620, -0.1923390, 0.1497640, 0.1792778, 0.1424335, -0.1931533, 0.1366939, 0.2007806, 0.2218272, -0.1268131, 0.2373037, 0.0212715, -0.2701837, -0.1922885, -0.0350652, 0.2434472, -0.1147770, -0.0435152, -0.1694131, -0.0205323, 0.0273878, 0.0035079, -0.0274193, 0.0911281, 0.1254953, -0.0251459, 0.2229911, 0.0872305, 0.1199639, 0.2197553, -0.1916868, -0.0770025, -0.1409274, 0.1261752, 0.2264333, -0.0465369, 0.0076258, 0.1262752, 0.1952620, -0.0224987, 0.1881456, -0.0363900, 0.1996294, -0.0478531, 0.0620196))
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s49,
    done => done_s50,
    start => start_s51,
    ack => ack_s52,
    in_a => in_a_s53,
    out_a => out_a_s54,
    out_offset => out_offset_s55,
    simd_offset => simd_offset_s56,
    op_argument => op_argument_s57,
    op_result => op_result_s58,
    op_send => op_send_s59,
    op_receive => op_receive_s60
);
conv_to_fc_interlayer_u138 : conv_to_fc_interlayer generic map(
    channels => 10,
    channel_width => 8,
    layer_size => 7,
    fc_simd => 70
) port map(
    clk => clk,
    ready => ready_s139,
    done => done_s140,
    start => start_s141,
    ack => ack_s142,
    din => din_s143,
    dout => dout_s144,
    wr_addr => wr_addr_s145,
    rd_addr => rd_addr_s146,
    wren_in => wren_in_s147
);
bias_op_u61 : bias_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 13, frac => 15)),
    bias_spec => fixed_spec(fixed_spec'(int => 1, frac => 11)),
    biases => reals(reals'( -0.4303576, -0.3637567, -0.3914840, -0.4656740, -0.3534780, -0.2577450, -0.7783858, -0.3849082, -0.3757767, -0.4386353, -0.3143329, -0.6888475, -0.2492339, -0.4169823, -0.1258507, 0.0593796, -0.3067093, -0.7916161, -0.5134744, -0.5892171, -0.3995129, -0.2564527, -0.4102712, -0.6959279, -0.5062674, -0.4237090, -0.5224990, -0.3688354, -0.4979883, -0.2034408, -0.0357736, -0.7220469, -0.2233848, -0.3427513, -0.8202428, -0.4750255, -0.4662284, -0.5145087, -0.2851815, -0.6549429))
) port map(
    input => input_s62,
    offset => offset_s63,
    output => output_s64,
    op_send => op_send_s65,
    op_receive => op_receive_s66
);
relu_op_u67 : relu_op generic map(
    spec => fixed_spec(fixed_spec'(int => 14, frac => 15))
) port map(
    input => input_s68,
    output => output_s69,
    op_send => op_send_s70,
    op_receive => op_receive_s71
);
fc_layer_u72 : fc_layer generic map(
    input_width => 40,
    output_width => 10,
    simd_width => 10,
    input_spec => fixed_spec(fixed_spec'(int => 3, frac => 8)),
    weight_spec => fixed_spec(fixed_spec'(int => 2, frac => 6)),
    op_arg_spec => fixed_spec(fixed_spec'(int => 13, frac => 14)),
    output_spec => fixed_spec(fixed_spec'(int => 4, frac => 8)),
    n_weights => 400,
    pick_from_ram => false,
    weights_filename => "whatever",
    weight_values => reals(reals'( -0.8604600, 0.0463802, -0.9526252, 0.2115245, -1.1042989, 0.2500386, 0.2449825, -1.2655805, -0.0356142, -0.7283774, -1.1949919, 0.1654240, -0.7354884, -0.6740655, 0.0426578, -0.8763394, -1.0828230, 0.2296938, -0.8801801, 0.1629041, -0.4766511, -1.1921548, -1.3634456, -0.8700417, -0.1489989, 0.4128420, 0.5061616, -1.0217036, -0.2737932, 0.4142204, -0.5062813, 0.1920487, 0.1446232, -0.9703508, 0.1719468, -0.4527321, 0.2040390, -0.6192911, -0.5547584, -0.7857679, -0.9092683, -1.0261070, -1.0518352, 0.1917799, -1.1540393, 0.2546712, 0.2818768, -1.3327903, 0.1774581, -0.4995609, 0.3388270, -1.1481732, -0.4449528, -1.1219537, 0.3588556, -1.1836098, -0.6963025, -0.6518287, -0.0038507, 0.2785923, -0.8182174, 0.0840578, 0.1417176, 0.1732988, -1.1410141, 0.1362479, -1.0513281, 0.1754692, -0.9613819, -0.5428103, 0.6282824, 0.4265591, -0.8592541, -1.1281902, -1.1307584, -0.7719007, -0.7308800, 0.4381461, -0.9756523, -0.6488369, 0.1509024, -1.1696488, -1.4116796, -1.1306336, -0.8685537, 0.0829138, 0.1709682, -0.9861229, -0.0672631, -1.0273036, 0.0412073, -0.6794091, 0.0620647, 0.0411900, -1.4078937, -0.8404651, -1.4215115, 0.0123338, -0.0456351, -0.7629471, -1.0308586, 0.2693282, -0.9134704, -1.1299140, 0.3381674, 0.2265147, -0.4619581, -0.5631486, 0.2162205, 0.2513451, -1.0674671, -0.5154473, -0.5848554, 0.1234185, 0.1370029, 0.1532462, -1.2637327, 0.1669483, -0.3473806, 0.1509154, -0.9451657, 0.4273389, -0.5616114, -0.9707852, -0.6142341, -0.8810729, -0.7353680, 0.4421622, -0.7914838, -0.5495354, -1.3439229, -0.9360925, -0.8824150, 0.2179996, 0.1320648, 0.2625083, -0.7462891, 0.2472340, 0.2184164, -0.5834519, 0.2898844, 0.1378301, -1.0320808, -1.5583655, -0.7843871, -0.6042159, 0.2990203, -0.9514294, 0.1331401, -1.3087777, -1.0304934, 0.5520027, -1.1480901, -1.3567516, -0.2893062, -1.1269530, -0.9875938, -0.7145211, 0.5733047, 0.4060538, -0.6350263, -1.1993052, -1.7174664, -1.0314001, -0.8426535, 0.2147859, 0.2769101, -1.2473031, 0.1642632, 0.0456816, 0.1695030, 0.1173766, 0.1105470, 0.0797785, -0.7650485, 0.1416692, 0.1631418, -0.6790126, -0.6570328, -0.7962485, -1.1881883, -0.6031290, -0.6913013, -0.5142890, 0.3187979, -0.7909168, -0.9549592, 0.2812263, -0.5949302, 0.2460957, -0.9187449, -0.6193160, 0.1640218, 0.1383213, -0.9331836, -0.9385080, -1.9472352, 0.1669588, 0.0162749, 0.0905766, -0.6559857, -1.2425879, -1.0069364, 0.2067174, 0.1591531, 0.1649268, -1.2618426, -0.6326240, 0.1457995, 0.1729100, -1.0007850, -0.9288440, 0.3379541, -0.3874722, -1.3610041, 0.2772114, -0.2059029, -0.8490391, 0.2711628, -0.6908261, 0.2250821, -0.9590064, 0.0717992, -0.9642665, -0.7023931, -0.4420470, 0.2429661, -1.2345413, 0.0236939, -1.1764069, -0.8260307, 0.1693618, 0.1668360, 0.0836271, 0.1392652, -0.8098346, -0.0867873, 0.1120075, -0.8099957, -0.8490582, -0.9422650, 0.1776808, 0.1622553, -0.7048568, 0.1993037, -1.0187081, -0.7643000, 0.1697624, 0.0149675, -0.7668450, -0.0900066, 0.1309751, -0.9010152, 0.1484603, -1.3679528, 0.1518742, -0.9994965, -0.7419205, -1.2232959, -0.4471471, -0.9069682, -0.2284389, 0.1666114, 0.1962885, -1.1407404, 0.1092049, -1.1328281, 0.1721341, 0.0711699, -0.6032202, -1.3022819, 0.1824711, -0.8252159, -0.4337380, -0.6271302, -0.7128643, -1.2357547, 0.3339511, -0.8253779, 0.1684327, -1.2951218, 0.3201509, -0.6163955, 0.2538179, 0.3384596, 0.2945586, -0.6828677, -0.4894696, -0.6898976, 0.1675055, -0.9637379, 0.1729572, 0.2076812, 0.1642146, 0.1962852, -0.9290428, -0.9730872, -0.2830532, 0.0929738, -0.7097578, -0.8830505, -1.4866589, -0.7905290, 0.5263599, -1.0412620, -0.7245772, -1.7259952, -0.8718196, 0.5189202, 0.4204054, 0.2140926, -0.9372647, -0.5365253, -0.9049960, 0.2038888, 0.1414681, -0.4307157, 0.1840671, -0.9900571, 0.1647475, 0.3848175, -0.8037407, 0.3507108, -0.5529093, -0.9784968, -0.9810251, -0.9555941, -0.6794043, 0.2657704, -0.8585753, -0.6444212, 0.0589940, 0.0866340, -1.2356504, 0.1557317, -0.6993470, 0.1942464, -0.7089474, 0.0571829, -0.7958655, -0.6335117, -0.5841568, 0.1501451, 0.0985995, 0.2071887, -0.7350762, 0.2350585, 0.1978747, -0.9323540, -0.8211558, -1.0994076, -0.9564958, 0.2297916, 0.2085882, -0.7832779, 0.1874181, -1.1850089, -0.5778830, -1.0604903, 0.2173264, 0.1446208, -1.3044430, -0.8866290, -1.4732434, 0.1168055, -0.0258223, 0.2029440, -0.7261818, -0.8072184, -0.7666973, -0.4496007, 0.1270381, 0.0905949, -1.0138381, 0.1550478, -0.4822470, 0.1790110, -0.6260436, -0.7401367, -0.6430855, 0.5318609, -1.5003012, -0.3445090, 0.4537367, -0.5354945, -0.8754864, -1.2943360, -0.7232026, -0.8294089, 0.4065037, 0.2561508, -0.8657771, 0.2078299, -0.4730174, -0.7934895, -0.9461973, -0.6789944, 0.2397927, -0.8740532, 0.0702637))
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s73,
    done => done_s74,
    start => start_s75,
    ack => ack_s76,
    in_a => in_a_s77,
    out_a => out_a_s78,
    out_offset => out_offset_s79,
    simd_offset => simd_offset_s80,
    op_argument => op_argument_s81,
    op_result => op_result_s82,
    op_send => op_send_s83,
    op_receive => op_receive_s84
);
fc_to_fc_interlayer_u149 : fc_to_fc_interlayer generic map(
    width => 40,
    word_size => 11
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s150,
    done => done_s151,
    start => start_s152,
    ack => ack_s153,
    previous_a => previous_a_s154,
    next_a => next_a_s155
);
bias_op_u85 : bias_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 13, frac => 14)),
    bias_spec => fixed_spec(fixed_spec'(int => 1, frac => 11)),
    biases => reals(reals'( 0.8162096, -0.2501919, -0.3209949, -0.5684234, -0.3526796, -0.8672848, 0.0149040, -0.4194804, 0.4514914, 0.5552633))
) port map(
    input => input_s86,
    offset => offset_s87,
    output => output_s88,
    op_send => op_send_s89,
    op_receive => op_receive_s90
);
sigmoid_op_u91 : sigmoid_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 14, frac => 14)),
    output_spec => fixed_spec(fixed_spec'(int => 4, frac => 8)),
    step_precision => 2,
    bit_precision => 16
) port map(
    clk => clk,
    input => input_s92,
    output => output_s93,
    op_send => op_send_s94,
    op_receive => op_receive_s95
);

din_s111 <= dout_s7;
ack_s4 <= load_done_s17;
done_s109 <= done_s2;
ready_s98 <= ready_s1;
rd_addr_s104 <= addr_s8;
start_s3 <= start_s100;
din_s6 <= dout_s102;
row_s115 <= row_s10;
wren_s116 <= wren_s11;
wr_addr_s113 <= out_addr_s9;
din_s121 <= dout_s19;
ack_s16 <= load_done_s29;
done_s119 <= done_s14;
ready_s108 <= ready_s13;
rd_addr_s114 <= addr_s20;
start_s15 <= start_s110;
din_s18 <= dout_s112;
row_s125 <= row_s22;
wren_s126 <= wren_s23;
wr_addr_s123 <= out_addr_s21;
din_s131 <= dout_s31;
ack_s28 <= load_done_s41;
done_s129 <= done_s26;
ready_s118 <= ready_s25;
rd_addr_s124 <= addr_s32;
start_s27 <= start_s120;
din_s30 <= dout_s122;
row_s135 <= row_s34;
wren_s136 <= wren_s35;
wr_addr_s133 <= out_addr_s33;
din_s143 <= dout_s43;
ack_s40 <= ack_s142;
done_s140 <= done_s38;
ready_s128 <= ready_s37;
rd_addr_s134 <= addr_s44;
start_s39 <= start_s130;
din_s42 <= dout_s132;
wren_in_s147 <= wren_s47;
wr_addr_s145 <= out_addr_s45;
previous_a_s154 <= out_a_s54;
ack_s52 <= ack_s153;
done_s151 <= done_s50;
in_a_s53 <= dout_s144;
start_s51 <= start_s141;
ready_s139 <= ready_s49;
rd_addr_s146 <= std_logic_vector(resize(unsigned(simd_offset_s56), rd_addr_s146'length));
input_s62 <= op_argument_s57;
op_receive_s66 <= op_send_s59;
op_receive_s60 <= op_send_s70;
input_s68 <= output_s64;
op_receive_s71 <= op_send_s65;
offset_s63 <= out_offset_s55;
op_result_s58 <= resize(output_s69, mk(fixed_spec(fixed_spec'(int => 3, frac => 8))));
in_a_s77 <= next_a_s155;
start_s75 <= start_s152;
ready_s150 <= ready_s73;
input_s86 <= op_argument_s81;
op_receive_s90 <= op_send_s83;
op_receive_s84 <= op_send_s94;
input_s92 <= output_s88;
op_receive_s95 <= op_send_s89;
offset_s87 <= out_offset_s79;
op_result_s82 <= resize(output_s93, mk(fixed_spec(fixed_spec'(int => 4, frac => 8))));

done_s99 <= start;
out_a <= out_a_s78;
end system;
